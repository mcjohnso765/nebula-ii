* NGSPICE file created from team_03_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

.subckt team_03_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ ncs vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08326__A3 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06883_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] team_03_WB.instance_to_wrap.core.decoder.inst\[27\]
+ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__or3_1
X_09671_ _05089_ _05091_ _05095_ _05098_ net556 net566 vssd1 vssd1 vccd1 vccd1 _05613_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11866__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08731__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ _04558_ _04563_ net870 vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13840__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11881__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__B _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11618__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ net850 _04493_ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07298__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _03443_ _03445_ net803 vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__o21a_1
X_08484_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07435_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\] net756
+ net725 _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1071_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout427_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13350__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08247__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\]
+ net757 vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09105_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\] net932
+ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07297_ net1158 _03237_ _03238_ _03234_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__o22a_1
XANTENNA__14346__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09974__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09036_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\]
+ net981 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11149__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout796_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold340 team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\] vssd1
+ vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold351 team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\] vssd1
+ vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06899__A _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold362 team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\] vssd1
+ vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07494__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold373 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\] vssd1
+ vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _02618_ vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__A2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\] vssd1
+ vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 _02846_ vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07773__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08970__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 net832 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_4
X_09938_ _05873_ net1793 net293 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
Xfanout842 _06303_ vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout853 net854 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__clkbuf_4
Xfanout864 net866 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__clkbuf_8
Xfanout875 net884 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_2
XANTENNA__11029__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__B1 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout886 net887 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__buf_2
Xfanout897 net900 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_2
X_09869_ net582 _05597_ _05804_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_99_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1040 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\] vssd1
+ vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\] vssd1
+ vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\] vssd1
+ vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net638 _06709_ net479 net380 net2329 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12880_ net1428 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
Xhold1073 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\] vssd1
+ vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\] vssd1
+ vssd1 vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\] vssd1
+ vssd1 vccd1 vccd1 net2679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11831_ net648 _06666_ net459 net328 net1817 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07289__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ clknet_leaf_85_wb_clk_i _02314_ _00915_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11762_ _06590_ net461 net340 net2334 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13501_ net1323 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] _05518_ net600 vssd1
+ vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14481_ clknet_leaf_94_wb_clk_i _02245_ _00846_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\]
+ sky130_fd_sc_hd__dfrtp_1
X_11693_ _06735_ net390 net346 net2526 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input92_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ net1425 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XANTENNA__12034__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10644_ net1203 net2675 net839 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08354__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13363_ net1332 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
X_10575_ net1928 net534 net595 _05885_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ net1483 vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_2
XFILLER_0_49_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15064__1445 vssd1 vssd1 vccd1 vccd1 _15064__1445/HI net1445 sky130_fd_sc_hd__conb_1
XANTENNA__07461__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ net1371 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13294_ net1392 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15033_ clknet_leaf_33_wb_clk_i _02753_ _01398_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11919__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12245_ net1751 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09753__A2 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ net1706 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08961__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ net625 _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__nor2_1
XANTENNA__06972__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11848__A0 _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ net515 net658 _06606_ net427 net2611 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07516__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11654__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _02888_ net1991 net288 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__mux2_1
XANTENNA__10520__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14817_ clknet_leaf_31_wb_clk_i net1775 _01182_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08477__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14748_ clknet_leaf_116_wb_clk_i _02512_ _01113_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14679_ clknet_leaf_52_wb_clk_i _02443_ _01044_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06991__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07220_ _03160_ _03161_ net1151 vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__o21a_1
XANTENNA__12025__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08229__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07151_ net1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\]
+ net879 _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ net611 _03023_ _02995_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11551__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07984_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\]
+ net900 vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_1475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09723_ _03759_ _04893_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__nor2_1
X_06935_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\]
+ net769 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__mux2_1
XANTENNA__11839__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_A net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13345__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ net592 _05584_ _05585_ _05595_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__o31a_2
XANTENNA__10511__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\] _02794_ _02806_
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__and3_4
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08605_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\]
+ net973 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
X_09585_ _05420_ _05525_ net570 vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout544_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1286_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08536_ net545 _04476_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08468__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10814__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[27\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout711_A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout809_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12016__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07418_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\]
+ net886 net1116 vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08398_ _04334_ _04339_ net871 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
XANTENNA__07691__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\] net1115
+ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o221a_1
XANTENNA__10578__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ _06092_ _06187_ _06101_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_27_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07994__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09019_ _04959_ _04960_ net862 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10291_ _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__or2_1
XANTENNA__10643__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _06771_ net482 net368 net2601 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\] vssd1
+ vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\] vssd1
+ vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\] vssd1
+ vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07746__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout650 _06457_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
Xfanout661 net662 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_4
Xfanout672 net673 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_4
X_13981_ clknet_leaf_66_wb_clk_i _01745_ _00346_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09499__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout694 _06562_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_8
X_12932_ net1311 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XANTENNA__08349__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12863_ net1378 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14602_ clknet_leaf_2_wb_clk_i _02366_ _00967_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11058__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11814_ _06642_ net473 net330 net1901 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__a22o_1
X_12794_ net1371 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14533_ clknet_leaf_108_wb_clk_i _02297_ _00898_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11745_ _06566_ net456 net337 net2304 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464_ clknet_leaf_132_wb_clk_i _02228_ _00829_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ net1038 net694 _06803_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13415_ net1424 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10627_ net1611 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] net835 vssd1 vssd1 vccd1
+ vccd1 _02501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10569__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14395_ clknet_leaf_28_wb_clk_i _02159_ _00760_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ net1291 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
X_10558_ net2037 net534 net595 _05868_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11649__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ net1396 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
X_10489_ net111 net1025 net905 net1802 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15016_ clknet_leaf_62_wb_clk_i _02736_ _01381_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09119__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ net1694 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11533__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ net1624 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07832__S1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14041__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08698__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11836__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_133_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09370_ _04071_ _05159_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15179__1560 vssd1 vssd1 vccd1 vccd1 _15179__1560/HI net1560 sky130_fd_sc_hd__conb_1
X_08321_ net944 _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\]
+ net946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\] net913
+ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07673__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07203_ net801 _03143_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\]
+ net947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\] net913
+ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12013__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__S0 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07134_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\]
+ net779 net1126 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07425__B1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06941__S net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11772__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07065_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\]
+ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput220 net220 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_101_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput231 net231 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput242 net242 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_100_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput253 net253 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__A1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout494_A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08925__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1201_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout661_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09025__S0 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ net745 _03905_ _03906_ _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09706_ _05211_ _05276_ _05209_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a21oi_1
X_06918_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\] net730
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07898_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\] net781
+ _03839_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__a21o_1
XANTENNA__08153__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ _05406_ _05408_ net555 vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__mux2_1
X_15063__1444 vssd1 vssd1 vccd1 vccd1 _15063__1444/HI net1444 sky130_fd_sc_hd__conb_1
X_06849_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] vssd1 vssd1 vccd1 vccd1
+ _02792_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout926_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09568_ _03904_ _04235_ _05509_ _02945_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09102__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08519_ net864 _04460_ _04455_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10638__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ net574 _05440_ _05439_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09653__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ net2404 net489 _06783_ net518 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08861__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11461_ net642 _06586_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ net1430 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_10412_ _05925_ _05945_ _06234_ _06235_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a22o_1
X_11392_ net509 net632 _06748_ net407 net2454 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a32o_1
X_14180_ clknet_leaf_12_wb_clk_i _01944_ _00545_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07967__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11763__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ net1254 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
X_10343_ _06148_ _06149_ _06178_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10971__A0 _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09169__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input55_A gpio_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ net1426 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
X_10274_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__inv_2
XANTENNA__14064__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07719__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net621 _06572_ net464 net365 net2160 vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__a32o_1
Xfanout1401 net1404 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__buf_4
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1412 net1432 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1423 net1425 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08392__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout480 net484 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 _06680_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13964_ clknet_leaf_9_wb_clk_i _01728_ _00329_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12915_ net1265 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
X_13895_ clknet_leaf_69_wb_clk_i _01659_ _00260_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13901__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11932__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ net1336 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07104__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ net1252 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14516_ clknet_leaf_92_wb_clk_i _02280_ _00881_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ net1961 _06491_ net341 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11451__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ clknet_leaf_99_wb_clk_i _02211_ _00812_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11659_ net2130 _06622_ net350 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07407__B1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14378_ clknet_leaf_4_wb_clk_i _02142_ _00743_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold906 team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\] vssd1
+ vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold917 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\] vssd1
+ vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold928 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\] vssd1
+ vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__B1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ net1318 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09698__A2_N _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold939 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\] vssd1
+ vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07422__A3 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10962__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _04809_ _04810_ _04770_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14557__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07821_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\] net760
+ net742 _03762_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07752_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\]
+ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__or2_1
XANTENNA__12003__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07683_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__and3_1
XANTENNA__10031__B net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13623__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _04816_ _05343_ _05361_ _05362_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06936__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09635__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\]
+ net983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\] net1071
+ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__o221a_1
XANTENNA__11143__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07646__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08843__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09284_ _04922_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08235_ net849 _04170_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout1151_A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08166_ net1220 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\]
+ net949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\] net930
+ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07949__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11745__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07117_ net722 _03058_ _03043_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__o21a_2
XFILLER_0_113_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08097_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\] net739
+ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__o221a_1
XFILLER_0_109_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09982__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07048_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _02808_ _02818_ net1138
+ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_100_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09020__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09166__A3 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10921__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08374__A1 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08999_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\]
+ net954 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08126__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[2\] net307 vssd1 vssd1
+ vccd1 vccd1 _06542_ sky130_fd_sc_hd__and2_1
XANTENNA__07234__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net1346 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10484__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__B1 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ clknet_leaf_83_wb_clk_i _01444_ _00045_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10892_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[15\] _05865_ net321 _06403_
+ net687 vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__a41o_1
XFILLER_0_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12631_ net1413 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XANTENNA__09087__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07637__B1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12562_ net1405 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ clknet_leaf_76_wb_clk_i _02065_ _00666_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11513_ _06629_ net2708 net395 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__mux2_1
X_12493_ net1301 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ clknet_leaf_9_wb_clk_i _01996_ _00597_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11444_ net2676 net399 _06761_ net518 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11199__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11736__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ clknet_leaf_113_wb_clk_i _01927_ _00528_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\]
+ sky130_fd_sc_hd__dfrtp_1
X_11375_ net1241 net831 net270 net666 vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10944__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ net1365 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
X_10326_ _06164_ _06165_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] net675
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ clknet_leaf_70_wb_clk_i _01858_ _00459_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11927__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ net1267 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09905__B _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ _04324_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] net671 vssd1
+ vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1220 net1223 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07706__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1231 net1233 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10188_ _03460_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1242 net1244 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
Xfanout1253 net1255 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__buf_4
XANTENNA__06915__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1264 net1266 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_4
Xfanout1275 net1276 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1286 net1295 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1297 net1317 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__buf_4
X_14996_ clknet_leaf_107_wb_clk_i net44 _01361_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08117__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13947_ clknet_leaf_28_wb_clk_i _01711_ _00312_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07325__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09865__B2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11662__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07876__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__D_N _05611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__A1 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ clknet_leaf_82_wb_clk_i _01642_ _00243_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10786__B net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ net1372 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08971__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07587__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ net1130 _03956_ _03960_ _03961_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold703 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\] vssd1
+ vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold714 team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\] vssd1
+ vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08053__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold725 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\] vssd1
+ vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
X_15062__1443 vssd1 vssd1 vccd1 vccd1 _15062__1443/HI net1443 sky130_fd_sc_hd__conb_1
XFILLER_0_106_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold736 team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\] vssd1
+ vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\] vssd1
+ vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\] vssd1
+ vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _03205_ net661 vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nor2_1
Xhold769 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07319__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13947__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\] net977
+ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or2_1
XANTENNA__09148__A3 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08356__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__B2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\] net943
+ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a221o_1
XANTENNA__11360__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07804_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\] net730
+ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a221o_1
XANTENNA__11138__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08784_ _04724_ _04725_ net864 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08108__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ net1139 _03672_ _03674_ _03676_ _02864_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a41o_1
XANTENNA__11112__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__S1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout457_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07867__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ net1166 team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\]
+ net885 net1115 vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09405_ _05164_ _05340_ _05345_ net582 vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o31a_1
X_07597_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout624_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1366_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09977__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09336_ _05235_ _05275_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__a21o_2
XFILLER_0_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ _05207_ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14722__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\]
+ net957 net1069 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux4_1
XANTENNA__09278__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ net567 _05134_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout993_A _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08149_ net930 _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10926__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11160_ net657 _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07229__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14872__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _04807_ net659 vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11091_ net830 net272 vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10651__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158__1539 vssd1 vssd1 vccd1 vccd1 _15158__1539/HI net1539 sky130_fd_sc_hd__conb_1
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08347__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ net15 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1
+ vccd1 vccd1 _02689_ sky130_fd_sc_hd__a22o_1
Xhold30 team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\] vssd1
+ vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\] vssd1
+ vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14850_ clknet_leaf_52_wb_clk_i net1882 _01215_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
Xhold52 team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\] vssd1
+ vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\] vssd1
+ vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold74 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\] vssd1
+ vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\] vssd1
+ vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ clknet_leaf_77_wb_clk_i _01565_ _00166_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold96 team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\] vssd1
+ vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ clknet_leaf_31_wb_clk_i _02545_ _01146_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net299 net2622 net449 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__mux2_1
XANTENNA__10887__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13732_ clknet_leaf_8_wb_clk_i _01496_ _00097_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07858__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ net512 net593 net265 net522 net1821 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a32o_1
XANTENNA__07322__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14252__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13663_ clknet_leaf_120_wb_clk_i _01427_ _00028_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10875_ net691 net318 net586 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_27_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12614_ net1419 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08807__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net1280 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07086__A1 net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12545_ net1287 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12476_ net1346 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XANTENNA__07200__S net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ clknet_leaf_65_wb_clk_i _01979_ _00580_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11427_ net633 net705 _06463_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__and3_4
XANTENNA__08035__B1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15195_ net1573 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10917__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__A _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ clknet_leaf_130_wb_clk_i _01910_ _00511_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09783__B1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11358_ net498 net615 _06731_ net405 net2519 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] _06150_ vssd1 vssd1
+ vccd1 vccd1 _06151_ sky130_fd_sc_hd__and2_1
X_14077_ clknet_leaf_66_wb_clk_i _01841_ _00442_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\]
+ sky130_fd_sc_hd__dfrtp_1
X_11289_ net1243 net834 _06536_ net669 vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__and4_2
XFILLER_0_67_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ net1314 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11342__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 _02791_ vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1061 net1063 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11893__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09550__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1083 net1085 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__buf_2
XANTENNA__08966__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10797__A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ clknet_leaf_31_wb_clk_i _02731_ _01344_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dfrtp_1
X_07520_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\] net1124
+ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a221o_1
XANTENNA__08510__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07451_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\]
+ net874 vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07382_ net808 _03319_ _03320_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__o22a_1
XANTENNA__11124__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10736__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08274__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09052_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\] net1074
+ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ net613 _03943_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__nor2_1
XANTENNA__14895__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08026__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\] vssd1
+ vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\] vssd1
+ vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\] vssd1
+ vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08577__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\] vssd1
+ vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold544 team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\] vssd1
+ vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11581__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold555 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\] vssd1
+ vssd1 vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold566 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\] vssd1
+ vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\] vssd1
+ vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\] vssd1
+ vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13348__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09954_ _05881_ net2015 net294 vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold599 team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\] vssd1
+ vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12252__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1114_A _02786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09037__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ _04841_ _04846_ net868 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09885_ _03137_ _04148_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nor2_1
Xhold1200 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\] vssd1
+ vssd1 vccd1 vccd1 net2784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1211 team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\] vssd1
+ vssd1 vccd1 vccd1 net2795 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ _02993_ net360 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nand2_2
Xhold1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\] vssd1
+ vssd1 vccd1 vccd1 net2806 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\] vssd1
+ vssd1 vccd1 vccd1 net2817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\] vssd1
+ vssd1 vccd1 vccd1 net2828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\] vssd1
+ vssd1 vccd1 vccd1 net2839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1 net2850
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1277 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1 net2861
+ sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ net1204 _04703_ _04705_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1288 team_03_WB.instance_to_wrap.core.pc.current_pc\[0\] vssd1 vssd1 vccd1 vccd1
+ net2872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ net817 _03651_ _03654_ _03659_ net717 vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_95_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08698_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\]
+ net978 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07649_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\]
+ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ net840 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ _04739_ _05258_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__nand2_1
XANTENNA__10646__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _06293_ _06300_ net1135 net1137 vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_88_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ net1250 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08017__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ net1287 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08568__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ clknet_leaf_81_wb_clk_i _01764_ _00365_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212_ net273 net2312 net490 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12192_ net1644 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08032__A3 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ net711 net694 net301 vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__or3b_1
XANTENNA__07240__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07256__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ net827 net278 vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__and2_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14618__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ net911 vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__inv_2
X_14902_ clknet_leaf_45_wb_clk_i _02665_ _01267_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14833_ clknet_leaf_31_wb_clk_i _02597_ _01198_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11627__A1 _06701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14768__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ clknet_4_6__leaf_wb_clk_i _02528_ _01129_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11976_ net280 net2728 net448 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15061__1442 vssd1 vssd1 vccd1 vccd1 _15061__1442/HI net1442 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13715_ clknet_leaf_113_wb_clk_i _01479_ _00080_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10927_ net690 _05718_ net587 vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__o21ai_1
X_14695_ clknet_leaf_43_wb_clk_i _02459_ _01060_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11940__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ clknet_leaf_71_wb_clk_i _01410_ _00011_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _06389_ _06390_ vssd1
+ vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__a21o_4
XFILLER_0_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08256__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13577_ net1397 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
X_10789_ _02932_ _06391_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__and2_4
XFILLER_0_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10063__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11241__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ net1427 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12459_ net1253 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08559__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11158__A3 _06656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__A _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ net1559 vssd1 vssd1 vccd1 vccd1 la_data_out[114] sky130_fd_sc_hd__buf_2
XFILLER_0_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09220__A2 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14129_ clknet_leaf_96_wb_clk_i _01893_ _00494_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07231__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout309 _06396_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07782__A2 _02821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11315__A0 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] net821 vssd1 vssd1 vccd1
+ vccd1 _02893_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07519__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09670_ _05187_ _05302_ _05305_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand3_1
X_06882_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] team_03_WB.instance_to_wrap.core.decoder.inst\[26\]
+ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1 vccd1 vccd1 _02824_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08731__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09381__A _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ net1064 _04561_ _04562_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08709__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\] net914
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__o221a_1
XFILLER_0_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07503_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\] net775
+ net750 _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o211a_1
XANTENNA__07298__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\]
+ net989 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11850__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07434_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\]
+ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15157__1538 vssd1 vssd1 vccd1 vccd1 _15157__1538/HI net1538 sky130_fd_sc_hd__conb_1
XFILLER_0_73_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07365_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\] net786
+ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout322_A net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A _02790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09104_ _05044_ _05045_ net850 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ net1149 _03235_ _03236_ net1112 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09035_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\]
+ net981 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1231_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11149__A3 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold330 team_03_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1 net1914
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold341 team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\] vssd1
+ vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold352 team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\] vssd1
+ vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__B net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\] vssd1
+ vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\] vssd1
+ vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold385 team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\] vssd1
+ vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\] vssd1
+ vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09990__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
Xfanout821 _02819_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08970__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _03563_ net661 vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nor2_1
Xfanout832 _06386_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__buf_4
XANTENNA__10109__A1 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout843 net844 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__buf_8
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 _04084_ vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_8
Xfanout865 net866 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13665__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ net359 _05107_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a21o_1
Xfanout887 net901 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__buf_4
Xhold1030 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\] vssd1
+ vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net900 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_8
Xhold1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\] vssd1
+ vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08819_ net1204 _04757_ _04758_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a31o_1
Xhold1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\] vssd1
+ vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1063 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\] vssd1
+ vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\] vssd1
+ vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09799_ _03489_ _04591_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__nand2_1
Xhold1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\] vssd1
+ vssd1 vccd1 vccd1 net2669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\] vssd1
+ vssd1 vccd1 vccd1 net2680 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ _06665_ net469 net329 net1889 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a22o_1
XANTENNA__10230__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07289__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11761_ net649 _06588_ net465 net340 net2114 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13500_ net1323 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_10712_ net1651 net531 net526 _06346_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08769__A1_N net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14480_ clknet_leaf_80_wb_clk_i _02244_ _00845_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\]
+ sky130_fd_sc_hd__dfrtp_1
X_11692_ _06734_ net392 net347 net2100 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08635__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13431_ net1421 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10643_ net1199 net2827 net840 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XANTENNA__12034__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08354__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input85_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ net1321 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ net1919 net537 net598 _05884_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15101_ net1482 vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_134_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ net1356 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07461__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ net1332 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ clknet_leaf_32_wb_clk_i _02752_ _01397_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__dfrtp_1
X_12244_ net1772 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12175_ net1615 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10405__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08961__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ net1242 net828 _06414_ net668 vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__or4_1
XANTENNA__07417__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06972__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09913__B _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ net1040 net834 _06545_ net669 vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08174__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _02921_ net1818 net291 vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14816_ clknet_leaf_56_wb_clk_i net1885 _01181_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08477__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ net619 _06736_ net458 net369 net1945 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a32o_1
X_14747_ clknet_leaf_14_wb_clk_i _02511_ _01112_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11670__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14678_ clknet_leaf_54_wb_clk_i _02442_ _01043_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13629_ net1404 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12025__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08229__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__A0 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__B1 _05907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07150_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\]
+ net1150 vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10587__B2 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__C1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07452__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07081_ net718 _03006_ _03015_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__o22a_4
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07204__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11000__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08401__B1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13688__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14933__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ net820 _03914_ _03924_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11845__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09722_ _05216_ _05662_ _05221_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13626__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ net818 _02875_ net723 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__a21o_1
XANTENNA__11839__A1 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__C1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B1 _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net359 _05587_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06865_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__or4bb_2
XANTENNA_fanout272_A _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\]
+ net973 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09584_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08535_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout537_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10275__A0 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08466_ net855 _04404_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10814__A2 _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07417_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08397_ net1215 _04337_ _04338_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout704_A _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10027__A0 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__A0 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09985__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07348_ net806 _03285_ _03286_ _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o22a_1
XANTENNA__10578__B2 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07279_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\] net732
+ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09018_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\] net981 net928
+ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a221o_1
XANTENNA__09286__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10290_ _05963_ _06128_ _06130_ net304 net305 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__a32o_1
XANTENNA__08190__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15060__1441 vssd1 vssd1 vccd1 vccd1 _15060__1441/HI net1441 sky130_fd_sc_hd__conb_1
Xhold160 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\] vssd1
+ vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 net235 vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07518__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\] vssd1
+ vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold193 team_03_WB.instance_to_wrap.CPU_DAT_I\[25\] vssd1 vssd1 vccd1 vccd1 net1777
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout640 net644 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_4
Xfanout662 _05860_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_4
X_13980_ clknet_leaf_120_wb_clk_i _01744_ _00345_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_2
XANTENNA__08156__C1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_4
Xfanout695 net700 vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__clkbuf_4
X_12931_ net1300 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07903__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06880__A_N _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12862_ net1414 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14601_ clknet_leaf_60_wb_clk_i _02365_ _00966_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\]
+ sky130_fd_sc_hd__dfstp_1
X_11813_ net648 _06640_ net460 net328 net1847 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a32o_1
XANTENNA__11058__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12793_ net1355 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XANTENNA__11490__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14532_ clknet_leaf_19_wb_clk_i _02296_ _00897_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\]
+ sky130_fd_sc_hd__dfrtp_1
X_11744_ _06565_ net471 net339 net2528 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07131__B1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08365__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ clknet_leaf_114_wb_clk_i _02227_ _00828_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\]
+ sky130_fd_sc_hd__dfrtp_1
X_11675_ net2436 _06633_ net350 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08306__S0 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ net1421 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ net1692 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] net835 vssd1 vssd1 vccd1
+ vccd1 _02502_ sky130_fd_sc_hd__mux2_1
X_14394_ clknet_leaf_21_wb_clk_i _02158_ _00759_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11766__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ net1292 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
X_10557_ net2852 net535 net596 _05861_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XANTENNA__12615__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09908__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13276_ net1395 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XANTENNA__11518__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ net112 net1025 net905 net1850 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15015_ clknet_leaf_38_wb_clk_i _02735_ _01380_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dfrtp_1
X_12227_ net1725 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07737__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net1688 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13980__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net265 net2697 net422 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15156__1537 vssd1 vssd1 vccd1 vccd1 _15156__1537/HI net1537 sky130_fd_sc_hd__conb_1
X_12089_ net634 _06656_ net472 net446 net1812 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07444__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08698__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07163__B _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08320_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08251_ _04187_ _04192_ net867 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__mux2_1
XANTENNA__11413__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A0 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__B1 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\] net737
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ net929 _04122_ _04123_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10029__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08848__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07133_ net1132 _03074_ net719 vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11221__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07619__A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ _02998_ _02999_ _03004_ _03005_ net1111 net1131 vssd1 vssd1 vccd1 vccd1 _03006_
+ sky130_fd_sc_hd__mux4_1
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11509__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput221 net221 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput232 net232 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
XFILLER_0_3_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput243 net243 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput254 net254 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1027_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10732__A1 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06985__D_N team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\]
+ net897 net1128 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a211o_1
XFILLER_0_96_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09025__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _05646_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__inv_2
X_06917_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\] net747
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11288__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\]
+ net880 _02870_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1396_A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ net571 _05486_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
X_06848_ net1232 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07361__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09567_ _03904_ _04235_ _04816_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout821_A _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__A0 _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout919_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08518_ _04456_ _04457_ _04459_ _04458_ net920 net859 vssd1 vssd1 vccd1 vccd1 _04460_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ _04448_ _04534_ net564 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08185__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09653__A2 _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__A0 _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08449_ net931 _04389_ _04390_ net850 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__o211a_1
XANTENNA__11460__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08861__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13853__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ net520 net634 _06585_ net400 net2192 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a32o_1
XFILLER_0_110_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11748__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ _06002_ _06004_ _06068_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08613__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ net1243 net833 _06545_ net667 vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__and4_1
XANTENNA__10654__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ net1248 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
X_10342_ team_03_WB.instance_to_wrap.core.pc.current_pc\[24\] _06148_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14209__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13061_ net1272 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
X_10273_ _04070_ _06113_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12012_ _06761_ net481 net367 net2511 vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a22o_1
Xfanout1402 net1404 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__buf_4
XANTENNA_input48_A gpio_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1413 net1415 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__buf_4
XANTENNA__11920__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1424 net1425 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_39_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout481 net484 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07264__A team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 _06680_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963_ clknet_leaf_17_wb_clk_i _01727_ _00328_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10487__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12914_ net1398 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
X_13894_ clknet_leaf_76_wb_clk_i _01658_ _00259_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12845_ net1290 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12776_ net1293 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07104__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11987__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ net2828 net300 net343 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14515_ clknet_leaf_115_wb_clk_i _02279_ _00880_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08852__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09919__A _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14446_ clknet_leaf_73_wb_clk_i _02210_ _00811_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\]
+ sky130_fd_sc_hd__dfrtp_1
X_11658_ net2108 _06479_ net351 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ net1710 team_03_WB.instance_to_wrap.CPU_DAT_O\[20\] net835 vssd1 vssd1 vccd1
+ vccd1 _02519_ sky130_fd_sc_hd__mux2_1
XANTENNA__07407__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ clknet_leaf_59_wb_clk_i _02141_ _00742_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11589_ _06473_ net2574 net452 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold907 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\] vssd1
+ vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold918 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\] vssd1
+ vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07439__A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13328_ net1292 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
Xhold929 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\] vssd1
+ vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10962__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13259_ net1272 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08907__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06918__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10714__B2 _06347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ net1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\]
+ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07591__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07751_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__or3_1
XANTENNA__07018__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07605__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10478__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07682_ net1106 _03622_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ net1017 net821 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1
+ vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11690__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08518__S0 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__A _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09352_ _04178_ _05292_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__nor2_2
XFILLER_0_118_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08209__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11978__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ _04241_ _04244_ net869 vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11143__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07646__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11442__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ _03243_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08843__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ net1077 _04175_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06952__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08165_ _04104_ _04105_ _04106_ net930 net1208 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout402_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1144_A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07116_ net818 _03049_ _03052_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08096_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\] net727
+ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__o221a_1
XFILLER_0_31_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07047_ net718 _02982_ _02988_ _02973_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1311_A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1409_A net1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14501__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08359__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout771_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__C1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net1209 _04939_ _04938_ net1201 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__o211a_1
XANTENNA__07084__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07949_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\]
+ net887 _03890_ net1145 vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10960_ net268 net2435 net522 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07334__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07885__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ net325 _05550_ _05560_ net326 _05557_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__a221o_1
XANTENNA__11681__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net317 _05846_ net320 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__o31a_1
XANTENNA__10649__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ net1345 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input102_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09087__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11969__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ net1312 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07637__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10641__A0 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14300_ clknet_leaf_128_wb_clk_i _02064_ _00665_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\]
+ sky130_fd_sc_hd__dfrtp_1
X_11512_ _06519_ net2387 net395 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12492_ net1296 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
X_15155__1536 vssd1 vssd1 vccd1 vccd1 _15155__1536/HI net1536 sky130_fd_sc_hd__conb_1
XANTENNA__14031__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14231_ clknet_leaf_75_wb_clk_i _01995_ _00596_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\]
+ sky130_fd_sc_hd__dfrtp_1
X_11443_ net656 _06570_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11197__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ clknet_leaf_104_wb_clk_i _01926_ _00527_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11736__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11374_ net508 net632 _06739_ net407 net1927 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10944__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08081__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ net1357 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10325_ net282 _06152_ _06161_ net675 vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__o31a_1
XANTENNA__07270__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14093_ clknet_leaf_106_wb_clk_i _01857_ _00458_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13044_ net1324 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
X_10256_ _06096_ _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__C _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1210 net1211 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1221 net1223 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1232 net1233 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_4
X_10187_ _04591_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] net672 vssd1
+ vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__mux2_1
Xfanout1243 net1244 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1254 net1255 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__buf_2
Xfanout1265 net1266 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
Xfanout1276 net1277 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
Xfanout1287 net1289 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
X_14995_ clknet_leaf_126_wb_clk_i net43 _01360_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1298 net1299 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__buf_4
XFILLER_0_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08748__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ clknet_leaf_7_wb_clk_i _01710_ _00311_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07325__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09865__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13877_ clknet_leaf_89_wb_clk_i _01641_ _00242_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10786__C net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12828_ net1341 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08825__B1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ net1417 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10632__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08553__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ clknet_leaf_60_wb_clk_i _02193_ _00794_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08589__C1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold704 team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\] vssd1
+ vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\] vssd1
+ vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold726 team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\] vssd1
+ vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\] vssd1
+ vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09970_ _05889_ net1922 net293 vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold748 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\] vssd1
+ vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\] vssd1
+ vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08921_ net439 net431 net588 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nor3_1
XFILLER_0_81_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09002__B1 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08852_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\] net925
+ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07564__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11360__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08761__C1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\] net747
+ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a221o_1
X_08783_ net1213 _04721_ _04722_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand3_1
XANTENNA__11138__B net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13634__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\] net789
+ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07316__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07867__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07665_ net1078 net885 team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\]
+ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout352_A _06805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15215__1579 vssd1 vssd1 vccd1 vccd1 _15215__1579/HI net1579 sky130_fd_sc_hd__conb_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _05164_ _05340_ _05345_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07596_ _03534_ _03537_ net819 vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09335_ _05204_ _05209_ _05213_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1359_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11966__A3 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _05041_ _05206_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08217_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\]
+ net973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09197_ net557 _05136_ _05138_ net573 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09993__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08148_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\] net949 net913
+ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout986_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07252__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08079_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\]
+ net890 _04020_ net1144 vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10110_ team_03_WB.instance_to_wrap.core.pc.current_pc\[0\] net659 vssd1 vssd1 vccd1
+ vccd1 _05954_ sky130_fd_sc_hd__nor2_1
X_11090_ _06479_ net2610 net423 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__S0 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net16 net1032 net906 net2282 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__o22a_1
XANTENNA__07555__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[10\] vssd1 vssd1 vccd1
+ vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold31 team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\] vssd1
+ vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold42 team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\] vssd1
+ vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\] vssd1
+ vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\] vssd1
+ vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\] vssd1
+ vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 net229 vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ clknet_leaf_18_wb_clk_i _01564_ _00165_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold97 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[14\] vssd1 vssd1 vccd1
+ vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ clknet_leaf_56_wb_clk_i _02544_ _01145_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11992_ net271 net2706 net448 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10887__B _05811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__A2 _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__C_N _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13731_ clknet_leaf_24_wb_clk_i _01495_ _00096_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\]
+ sky130_fd_sc_hd__dfrtp_1
X_10943_ net829 _06527_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13662_ clknet_leaf_77_wb_clk_i _01426_ _00027_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10874_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[18\] net308 net685 vssd1
+ vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ net1276 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08807__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13593_ net1281 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10614__A0 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08902__S0 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ net1379 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07086__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ net1360 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11426_ net296 net2437 net403 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__mux2_1
X_14214_ clknet_leaf_86_wb_clk_i _01978_ _00579_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\]
+ sky130_fd_sc_hd__dfrtp_1
X_15194_ net910 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10917__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14145_ clknet_leaf_0_wb_clk_i _01909_ _00510_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07243__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11938__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10842__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net710 _06468_ net695 vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__and3_1
XANTENNA__09916__B _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08820__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07794__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] _06148_ _06149_ vssd1
+ vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__and3_1
XANTENNA__07717__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__C1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ clknet_leaf_119_wb_clk_i _01840_ _00441_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\]
+ sky130_fd_sc_hd__dfrtp_1
X_11288_ net507 net630 _06711_ net416 net2270 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09535__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ net1267 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
X_10239_ _06004_ _06069_ _06077_ _06079_ _06075_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_98_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11342__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1040 _02793_ vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08743__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1051 net1053 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1073 net1076 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_4
XANTENNA__11673__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1084 net1085 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_2
Xfanout1095 net1098 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_2
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14978_ clknet_leaf_31_wb_clk_i _02730_ _01343_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10797__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13929_ clknet_leaf_58_wb_clk_i _01693_ _00294_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07450_ net1083 net889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10853__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07381_ net744 _03321_ _03322_ net805 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11124__D net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09120_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11948__A3 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08274__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\] net1207
+ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11140__C net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08026__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold501 team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\] vssd1
+ vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold512 team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\] vssd1
+ vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11848__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\] vssd1
+ vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13629__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold534 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\] vssd1
+ vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09774__B2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold545 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\] vssd1
+ vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 net204 vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold567 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\] vssd1
+ vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\] vssd1
+ vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _03984_ net661 vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__nor2_2
Xhold589 team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\] vssd1
+ vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ net1210 _04844_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__o21a_1
XANTENNA__06888__D _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _05283_ _05290_ _05599_ net583 vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout1107_A _02786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1201 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\] vssd1
+ vssd1 vccd1 vccd1 net2785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1212 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\] vssd1
+ vssd1 vccd1 vccd1 net2796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\] vssd1
+ vssd1 vccd1 vccd1 net2807 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ net585 _04775_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\] vssd1
+ vssd1 vccd1 vccd1 net2818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15154__1535 vssd1 vssd1 vccd1 vccd1 _15154__1535/HI net1535 sky130_fd_sc_hd__conb_1
Xhold1245 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\] vssd1
+ vssd1 vccd1 vccd1 net2829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11583__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1256 team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\] vssd1
+ vssd1 vccd1 vccd1 net2840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\] vssd1
+ vssd1 vccd1 vccd1 net2851 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ net1214 _04706_ _04707_ net1072 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__o211a_1
Xhold1278 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1 net2862
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1 net2873
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07362__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07717_ net813 _03656_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or3_1
XANTENNA__11636__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ net860 _04635_ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout734_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09988__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10844__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\]
+ net760 vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07579_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\] net798
+ _02869_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ _04808_ _04812_ _04811_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07068__A2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ team_03_WB.instance_to_wrap.core.i_hit _05914_ vssd1 vssd1 vccd1 vccd1 _06300_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07301__S _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ _04294_ _05189_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12260_ net1311 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11211_ _06468_ net2256 net490 vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13539__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ net1588 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07776__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11142_ net2308 net417 _06647_ net499 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a22o_1
XANTENNA__07537__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11059__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _06614_ net2548 net422 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ _05896_ _05897_ _05898_ _05901_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__or4_1
X_14901_ clknet_leaf_45_wb_clk_i _02664_ _01266_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11493__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08740__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14832_ clknet_leaf_62_wb_clk_i net1778 _01197_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_101_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11627__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14763_ clknet_leaf_16_wb_clk_i _02527_ _01128_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11975_ _06405_ net2855 net450 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13714_ clknet_leaf_100_wb_clk_i _01478_ _00079_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ net297 net2540 net523 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__mux2_1
X_14694_ clknet_leaf_53_wb_clk_i _02458_ _01059_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13937__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13645_ net1402 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
XANTENNA__10837__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ _06380_ _06389_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or2_4
XFILLER_0_73_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11522__A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13576_ net1310 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
X_10788_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[31\] team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[31\]
+ net308 vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__C _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12527_ net1388 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09927__A _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08831__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net1261 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11668__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ net274 net2805 net402 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
X_15177_ net1558 vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_2
X_12389_ net1275 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XANTENNA__07231__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ clknet_leaf_82_wb_clk_i _01892_ _00493_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06950_ net609 _02888_ _02890_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__o21ai_1
X_14059_ clknet_leaf_17_wb_clk_i _01823_ _00424_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08977__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07519__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07881__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08716__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06881_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _02823_ sky130_fd_sc_hd__and2_1
XANTENNA__11866__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ net1213 _04559_ _04560_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14712__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\] net931
+ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__o221a_1
XANTENNA__11618__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07502_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\]
+ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10826__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ net871 _04420_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or3_1
XANTENNA__08495__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07433_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\] net756
+ net738 _03374_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08247__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07364_ net1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\]
+ net885 net1142 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__o31a_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ net1220 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\] net930
+ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\]
+ net777 net1126 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ net944 _04974_ _04975_ net854 vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11578__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\] vssd1
+ vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 net231 vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1224_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\] vssd1
+ vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\] vssd1
+ vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold364 net232 vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\] vssd1
+ vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout800 _02850_ vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_8
Xhold386 team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\] vssd1
+ vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold397 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\] vssd1
+ vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _02848_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09936_ _05872_ net1796 net292 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__mux2_1
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_4
Xfanout833 net834 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_4
XANTENNA__06981__A1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout844 _04097_ vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__buf_8
XANTENNA__07791__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout855 net856 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_4
Xfanout866 _04082_ vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_8
X_09867_ net325 _05484_ _05495_ net327 _05808_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__a221o_1
XANTENNA__11857__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_A _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1020 team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\] vssd1
+ vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout888 net892 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_2
Xfanout899 net900 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1031 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\] vssd1
+ vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\] vssd1
+ vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\] vssd1
+ vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ net1216 _04756_ _04759_ net1072 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__o211a_1
Xhold1064 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\] vssd1
+ vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net581 _05739_ net359 vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__o21a_1
Xhold1075 team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\] vssd1
+ vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\] vssd1
+ vssd1 vccd1 vccd1 net2670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\] vssd1
+ vssd1 vccd1 vccd1 net2681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08749_ net1214 _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__and3_1
XANTENNA__10817__A0 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11760_ _06587_ net480 net338 net2439 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10711_ _02771_ _05499_ net600 vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07820__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ _06733_ net387 net345 net2386 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13430_ net1329 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
X_10642_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] team_03_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ net840 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XANTENNA__12034__A2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11061__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ net1288 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ net1974 net535 net596 _05883_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ net1481 vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_2
X_12312_ net1368 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13292_ net1332 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input78_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ clknet_leaf_41_wb_clk_i _02751_ _01396_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__dfrtp_1
X_12243_ net1758 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13269__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07749__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07267__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12174_ net1600 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ net2836 net417 _06637_ net496 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12901__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06972__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14735__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ net2317 net426 _06605_ net510 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09913__C _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _03488_ net2033 net289 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08098__A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10520__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14815_ clknet_leaf_62_wb_clk_i _02579_ _01180_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08477__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14746_ clknet_leaf_118_wb_clk_i _02510_ _01111_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11958_ net641 _06735_ net481 net371 net2048 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a32o_1
XANTENNA__09674__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07685__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ net298 net2524 net524 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__mux2_1
X_14677_ clknet_leaf_54_wb_clk_i _02441_ _01042_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11889_ net615 _06698_ net457 net377 net2094 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__a32o_1
XANTENNA__12348__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08229__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13628_ net1333 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11233__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07437__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13559_ net1404 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15153__1534 vssd1 vssd1 vccd1 vccd1 _15153__1534/HI net1534 sky130_fd_sc_hd__conb_1
X_07080_ net818 _03021_ net723 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__C_N net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07982_ net815 _03919_ _03921_ _03923_ net719 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__o41a_1
XFILLER_0_103_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12811__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06933_ net1110 _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__a21o_1
X_09721_ _05216_ _05221_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11427__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _05513_ _05545_ _05550_ net326 _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__a221o_1
X_06864_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10511__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08603_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\]
+ net974 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
X_09583_ net555 _05095_ _05524_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a21boi_2
XANTENNA__11146__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08534_ net437 net429 _04475_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__or3_4
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08468__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10985__B net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08465_ net850 _04405_ _04406_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout432_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1174_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11162__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08396_ net1062 _04335_ _04336_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07691__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10027__A1 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ net737 _03287_ _03288_ net801 vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10578__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__B1 _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07278_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\]
+ net778 vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ net944 _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11101__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11527__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07087__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\] vssd1
+ vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\] vssd1
+ vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\] vssd1
+ vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 net183 vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _02596_ vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07600__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 net633 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 net644 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_2
X_09919_ _03351_ net661 vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nor2_1
Xfanout652 _06457_ vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_4
Xfanout663 _04818_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
Xfanout674 _05948_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08156__B1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 net689 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11337__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout696 net700 vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__buf_2
X_12930_ net1353 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12861_ net1372 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
XANTENNA__09105__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14600_ clknet_leaf_34_wb_clk_i _02364_ _00965_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11812_ _06639_ net463 net331 net1864 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12792_ net1369 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XANTENNA__10895__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07550__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ clknet_leaf_25_wb_clk_i _02295_ _00896_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11463__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11743_ net1240 net701 _06803_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__or3_1
XANTENNA__07131__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11072__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14462_ clknet_leaf_57_wb_clk_i _02226_ _00827_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ net2253 _06632_ net349 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14288__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__A0 _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ net1329 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08306__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10625_ net1649 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] net835 vssd1 vssd1 vccd1
+ vccd1 _02503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14393_ clknet_leaf_93_wb_clk_i _02157_ _00758_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10569__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ team_03_WB.instance_to_wrap.core.ru.state\[5\] _06292_ net1137 vssd1 vssd1
+ vccd1 vccd1 _06299_ sky130_fd_sc_hd__and3b_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08631__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ net1289 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10487_ net2181 net1024 net905 net2031 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
X_13275_ net1396 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15014_ clknet_leaf_61_wb_clk_i _02734_ _01379_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12226_ net1663 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07428__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12157_ net1614 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _06629_ net2582 net422 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
X_12088_ _06788_ net465 net444 net2050 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__a22o_1
XANTENNA__08320__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ net496 net648 _06595_ net425 net2466 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a32o_1
XANTENNA__08698__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14729_ clknet_leaf_46_wb_clk_i _02493_ _01094_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11454__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08250_ net1208 _04190_ _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07201_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\] net724
+ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__o221a_1
XANTENNA__11206__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\] net948 net913
+ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11757__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07132_ net1112 _03068_ _03069_ _03070_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14900__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07976__A3 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07063_ _03000_ _03001_ net744 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
Xoutput211 net211 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput222 net222 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
Xoutput233 net233 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
Xoutput244 net244 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput255 net255 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11856__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10193__B1 _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07965_ net1099 net897 team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\]
+ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11157__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ net583 _05636_ _05637_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__a31o_2
XFILLER_0_78_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06916_ _02855_ _02857_ net803 vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07896_ _03835_ _03837_ net1112 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__a21o_1
XANTENNA__09886__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11693__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09635_ net570 _05487_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a21boi_1
X_06847_ net1215 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__inv_2
XANTENNA__10996__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07361__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09566_ _02992_ _04477_ _05125_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09061__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__A2 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ net568 net559 _04478_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout814_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08448_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\] net914
+ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _04317_ _04318_ _04320_ _04319_ net935 net857 vssd1 vssd1 vccd1 vccd1 _04321_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10410_ _06002_ _06004_ _06068_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14580__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ net511 net637 _06747_ net407 net2328 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10341_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] _06177_ net675 vssd1
+ vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13060_ net1316 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
X_10272_ _04070_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12011_ net617 _06569_ net456 net365 net2223 vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12451__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1403 net1404 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1414 net1415 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__buf_4
Xfanout1425 net1426 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08129__A0 _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout460 net485 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout471 net474 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07264__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 net484 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_4
Xfanout493 _06680_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ clknet_leaf_9_wb_clk_i _01726_ _00327_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09182__D _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12913_ net1312 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152__1533 vssd1 vssd1 vccd1 vccd1 _15152__1533/HI net1533 sky130_fd_sc_hd__conb_1
XANTENNA__11684__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13893_ clknet_leaf_108_wb_clk_i _01657_ _00258_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12844_ net1298 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12775_ net1399 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07104__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13678__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ clknet_leaf_101_wb_clk_i _02278_ _00879_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11726_ net2821 net272 net343 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14923__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14445_ clknet_leaf_106_wb_clk_i _02209_ _00810_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09919__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ net2817 _06621_ net348 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12626__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10608_ net1612 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] net838 vssd1 vssd1 vccd1
+ vccd1 _02520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ clknet_leaf_27_wb_clk_i _02140_ _00741_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11588_ _06468_ net2046 net452 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09801__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13327_ net1283 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
Xhold908 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\] vssd1
+ vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ net136 net1029 net1020 net1815 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
Xhold919 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\] vssd1
+ vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10146__A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10962__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13258_ net1248 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XANTENNA__08368__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12209_ net1620 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06918__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ net1271 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07040__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__A3 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07018__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _03688_ _03691_ net802 _03687_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14453__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\] net726
+ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07343__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09420_ _02782_ _02804_ net663 _05342_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08518__S1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _04178_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08302_ net853 _04242_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _03208_ _05146_ _02937_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08843__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11442__A3 _06569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08233_ net1212 _04174_ _04173_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10650__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10755__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11440__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10982__C net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08164_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08225__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10402__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ net809 _03054_ _03056_ net814 vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__o31a_1
XFILLER_0_113_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07949__A3 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _04034_ _04036_ net807 vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07803__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07046_ _02986_ _02987_ net818 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08359__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout597_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11586__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09020__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12271__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09056__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\]
+ net954 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
XANTENNA__07582__A1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07948_ net1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\]
+ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout931_A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ net723 _03806_ _03812_ _03820_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a22oi_4
XANTENNA__07334__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11130__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09618_ net565 _05469_ _05558_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a22o_1
XANTENNA__13820__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ net692 _05646_ net587 vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__o21a_1
XANTENNA__11418__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09087__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ _03529_ _04267_ net663 _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11969__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ net1427 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
XANTENNA__11053__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _06628_ net2689 net395 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ net1253 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ clknet_leaf_85_wb_clk_i _01994_ _00595_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11442_ net496 net617 _06569_ net397 net2292 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a32o_1
XANTENNA__11197__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14161_ clknet_leaf_96_wb_clk_i _01925_ _00526_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ net712 _06504_ net699 vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10944__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ _06162_ _06163_ net282 vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__a21bo_1
X_13112_ net1369 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XANTENNA_input60_A gpio_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14092_ clknet_leaf_8_wb_clk_i _01856_ _00457_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11496__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _03901_ _06095_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ net1264 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09011__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1 vccd1
+ vccd1 net1200 sky130_fd_sc_hd__buf_8
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ _06026_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1222 net1223 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07706__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1233 net1239 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__clkbuf_4
Xfanout1244 team_03_WB.instance_to_wrap.core.decoder.inst\[9\] vssd1 vssd1 vccd1 vccd1
+ net1244 sky130_fd_sc_hd__clkbuf_4
Xfanout1255 net1270 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_2
XFILLER_0_98_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1266 net1270 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__clkbuf_4
X_14994_ clknet_leaf_124_wb_clk_i net42 _01359_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1277 net1295 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_4
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_2
Xfanout1288 net1289 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_4
Xfanout1299 net1317 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08117__A3 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ clknet_leaf_111_wb_clk_i _01709_ _00310_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07325__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09865__A3 _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07876__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ clknet_leaf_90_wb_clk_i _01640_ _00241_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11409__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12827_ net1344 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12082__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ net1346 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08834__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10632__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11709_ _06459_ _06803_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ net1312 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06931__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14428_ clknet_leaf_127_wb_clk_i _02192_ _00793_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold705 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\] vssd1
+ vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
X_14359_ clknet_leaf_75_wb_clk_i _02123_ _00724_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08684__S0 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\] vssd1
+ vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\] vssd1
+ vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold738 team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\] vssd1
+ vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold749 team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\] vssd1
+ vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14819__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ net588 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08851_ _04791_ _04792_ net865 vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11896__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08761__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _03741_ _03743_ net803 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13843__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08782_ net1059 _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__nand2_1
XANTENNA__11138__C net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07913__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07733_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\] net763
+ net1011 vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07664_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09403_ _05343_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13993__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11154__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09069__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07595_ net804 _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__or3_1
XFILLER_0_88_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout345_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1087_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ _05235_ _05275_ _05213_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a21o_1
XANTENNA__08277__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11820__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09265_ _05041_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout512_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14349__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11170__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08216_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\]
+ net974 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__o221a_1
X_09196_ net548 _04771_ _05137_ net563 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08147_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15151__1532 vssd1 vssd1 vccd1 vccd1 _15151__1532/HI net1532 sky130_fd_sc_hd__conb_1
XFILLER_0_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07252__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\]
+ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ _02968_ _02970_ net746 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout979_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07095__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ net17 net1032 net906 net2047 vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08978__S1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\] vssd1
+ vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\] vssd1
+ vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\] vssd1
+ vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\] vssd1
+ vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold54 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\] vssd1
+ vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[4\] vssd1 vssd1 vccd1
+ vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold76 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\] vssd1
+ vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[16\] vssd1 vssd1 vccd1
+ vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11991_ _06487_ net2720 net451 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__mux2_1
Xhold98 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\] vssd1
+ vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ clknet_leaf_132_wb_clk_i _01494_ _00095_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10942_ _06524_ _06525_ _06526_ _06399_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__o211a_4
XFILLER_0_39_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ clknet_leaf_67_wb_clk_i _01425_ _00026_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[18\] net306 vssd1
+ vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ net1306 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12064__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08807__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13592_ net1263 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08902__S1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ net1374 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
XANTENNA__11811__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11080__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12474_ net1371 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13716__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ clknet_leaf_107_wb_clk_i _01977_ _00578_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\]
+ sky130_fd_sc_hd__dfrtp_1
X_11425_ net2864 net403 _06755_ net508 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a22o_1
X_15193_ net910 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10917__A2 _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ clknet_leaf_134_wb_clk_i _01908_ _00509_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07243__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ net495 net619 _06730_ net405 net1735 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09783__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08991__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and2_1
X_14075_ clknet_leaf_27_wb_clk_i _01839_ _00440_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11287_ net716 net269 net826 vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13026_ net1347 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
X_10238_ _03602_ _06073_ _06078_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__or3_1
XANTENNA__11878__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07546__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11342__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08743__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_4
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__clkbuf_4
X_10169_ _04893_ net673 vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1063 net1064 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_2
Xfanout1074 net1075 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08829__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1085 net1088 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__buf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_14977_ clknet_leaf_33_wb_clk_i _02729_ _01342_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11255__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13928_ clknet_leaf_35_wb_clk_i _01692_ _00293_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10853__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13859_ clknet_leaf_23_wb_clk_i _01623_ _00224_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12055__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07380_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\]
+ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10605__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09050_ net861 _04990_ _04991_ _04989_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__a31o_1
XANTENNA__07482__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08001_ net1212 _02821_ _03107_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14641__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__A2_N _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold502 team_03_WB.instance_to_wrap.core.ru.state\[3\] vssd1 vssd1 vccd1 vccd1 net2086
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold513 team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\] vssd1
+ vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07908__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\] vssd1
+ vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold535 team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\] vssd1
+ vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\] vssd1
+ vssd1 vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\] vssd1
+ vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold568 team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\] vssd1
+ vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09952_ _05880_ net1857 net295 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__mux2_1
Xhold579 team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\] vssd1
+ vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08903_ net1056 _04842_ _04843_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__or3_1
XANTENNA__11869__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _05283_ _05599_ _05290_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09082__S0 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11864__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1202 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\] vssd1
+ vssd1 vccd1 vccd1 net2786 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ net584 _02953_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__and2_1
Xhold1213 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\] vssd1
+ vssd1 vccd1 vccd1 net2797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10541__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\] vssd1
+ vssd1 vccd1 vccd1 net2808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1002_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\] vssd1
+ vssd1 vccd1 vccd1 net2819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11884__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1246 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\] vssd1
+ vssd1 vccd1 vccd1 net2830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14021__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1257 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\] vssd1
+ vssd1 vccd1 vccd1 net2841 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\] net1060
+ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a221o_1
Xhold1268 team_03_WB.instance_to_wrap.CPU_DAT_I\[31\] vssd1 vssd1 vccd1 vccd1 net2852
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout462_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1279 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\] vssd1
+ vssd1 vccd1 vccd1 net2863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11165__A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\] net789
+ net1037 _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__o211a_1
X_08696_ net852 _04636_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10844__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[21\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ net728 _03587_ _03588_ net1152 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_117_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1371_A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout727_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08474__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07578_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09317_ _04739_ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09462__A1 _05403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07473__B1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09248_ _04294_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08017__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09179_ net553 _04807_ net542 net583 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__o22a_1
XANTENNA__08648__S0 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13889__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07225__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _06453_ net2589 net490 vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__mux2_1
X_12190_ net1590 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11021__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07818__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08422__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09736__C net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08973__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11141_ net653 _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07029__S net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11072_ net830 net303 vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__and2_2
XANTENNA__11059__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput100 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_1
XANTENNA__07256__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ net91 net90 _05899_ _05900_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__or4_1
X_14900_ clknet_leaf_37_wb_clk_i _02663_ _01265_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__08725__B1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ clknet_leaf_62_wb_clk_i net1952 _01196_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14762_ clknet_leaf_42_wb_clk_i _02526_ _01127_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11974_ _06447_ _06751_ _06394_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__or3b_4
XFILLER_0_58_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13713_ clknet_leaf_96_wb_clk_i _01477_ _00078_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10835__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[23\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ net686 _06511_ _06512_ _06510_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__o31a_2
X_14693_ clknet_leaf_53_wb_clk_i _02457_ _01058_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07699__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13644_ net1310 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12037__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ _06380_ _06389_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11522__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13575_ net1424 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10787_ net315 net310 net319 vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__or3_1
XANTENNA__10063__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ net1340 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XANTENNA__11260__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ net1247 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11012__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ net301 net2832 net401 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__mux2_1
X_15176_ net1557 vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_2
X_12388_ net1303 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14127_ clknet_leaf_97_wb_clk_i _01891_ _00492_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ net1241 net831 net279 net666 vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09943__A _04029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ clknet_leaf_9_wb_clk_i _01822_ _00423_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07519__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ net1312 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XANTENNA__09662__B _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06880_ _02808_ _02817_ _02820_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\]
+ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__and4bb_1
XANTENNA__10523__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07463__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\]
+ net953 net914 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15150__1531 vssd1 vssd1 vccd1 vccd1 _15150__1531/HI net1531 sky130_fd_sc_hd__conb_1
XFILLER_0_37_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07501_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\] net794
+ net731 _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__o211a_1
X_08481_ _04421_ _04422_ net861 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__and3_1
XANTENNA__12028__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ net1138 _03297_ _03298_ net1152 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__o31a_1
XANTENNA__09444__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09102_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\] net995
+ net914 _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07455__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08798__A3 _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\]
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11859__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\] net928
+ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07638__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08404__C1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\] vssd1
+ vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 team_03_WB.instance_to_wrap.CPU_DAT_I\[6\] vssd1 vssd1 vccd1 vccd1 net1905
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold332 net209 vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\] vssd1
+ vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold354 team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\] vssd1
+ vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold365 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\] vssd1
+ vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\] vssd1
+ vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_A team_03_WB.instance_to_wrap.core.decoder.inst\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[24\] vssd1 vssd1 vccd1
+ vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold398 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\] vssd1
+ vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 _02849_ vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_8
X_09935_ _04069_ net660 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__nor2_2
XFILLER_0_99_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout812 _02847_ vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__clkbuf_8
Xfanout823 _06558_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10999__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout834 _06386_ vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_4
XANTENNA__11594__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06981__A2 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net849 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_8
Xfanout856 net858 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
XANTENNA__14537__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout867 net871 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__buf_4
X_09866_ _04824_ _05126_ _05371_ _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__a311o_1
XANTENNA__10514__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1010 team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\] vssd1
+ vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout878 net884 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1021 team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\] vssd1
+ vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08183__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout889 net892 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1032 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\] vssd1
+ vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\] net1060
+ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a221o_1
Xhold1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\] vssd1
+ vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _05110_ _05119_ _05130_ _05113_ net563 net572 vssd1 vssd1 vccd1 vccd1 _05739_
+ sky130_fd_sc_hd__mux4_1
Xhold1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\] vssd1
+ vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout844_A _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\] vssd1
+ vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07930__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\] vssd1
+ vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09999__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\] vssd1
+ vssd1 vccd1 vccd1 net2671 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\]
+ net975 net1072 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux4_1
Xhold1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\] vssd1
+ vssd1 vccd1 vccd1 net2682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08679_ net441 net433 _04620_ net553 vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__o31a_1
XANTENNA__10938__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10710_ net525 _06344_ _06345_ net530 net2345 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12019__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _06732_ net385 net344 net2014 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10641_ net1167 net1983 net839 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12034__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10045__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11061__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07446__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13360_ net1292 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
X_10572_ net1780 net537 net598 _05882_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a22o_1
XANTENNA__08643__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07997__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ net1414 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13291_ net1392 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15030_ clknet_leaf_54_wb_clk_i _02750_ _01395_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ net1756 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07548__A _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ net1673 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11124_ net280 net648 net703 net695 vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_1394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11055_ net654 net707 net268 net824 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__and4_1
XFILLER_0_99_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09913__D _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07283__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _03458_ net1705 net289 vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07921__A1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14814_ clknet_leaf_62_wb_clk_i net1762 _01179_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
X_14745_ clknet_leaf_13_wb_clk_i _02509_ _01110_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net634 _06734_ net472 net372 net2203 vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ net687 _06497_ _06498_ _06496_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__o31a_2
X_14676_ clknet_leaf_52_wb_clk_i _02440_ _01041_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ net617 _06697_ net456 net377 net2269 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a32o_1
XANTENNA__09774__A1_N net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13627_ net1313 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09426__A1 net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10839_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[22\] _05865_ net321 _06403_
+ net687 vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__a41o_1
XANTENNA__10149__A _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12025__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ net1424 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07988__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ net1375 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
X_13489_ net1334 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15159_ net1540 vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_0_11_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07981_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\] net798
+ _02871_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o211a_1
XANTENNA__13195__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _05217_ _05227_ _05660_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__and3_1
X_06932_ _02865_ _02866_ _02868_ net1123 net1156 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11839__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__B2 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09651_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11427__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06863_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\] vssd1 vssd1 vccd1
+ vccd1 _02805_ sky130_fd_sc_hd__nand3b_1
XANTENNA__07912__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ net921 _04542_ _04543_ net859 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ net550 _04417_ _05103_ net555 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a211o_1
XANTENNA__11146__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08533_ _04461_ _04474_ net843 vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__mux2_4
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09665__A1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\] net932
+ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11472__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10814__A4 _06403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11162__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07415_ net1080 net886 team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\]
+ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__o21a_1
XANTENNA__09417__A1 _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08395_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\]
+ net990 net1074 vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout425_A net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1167_A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07346_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\]
+ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11589__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07277_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\]
+ net777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\] net748
+ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1334_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\]
+ net981 vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11527__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold140 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\] vssd1
+ vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\] vssd1
+ vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\] vssd1
+ vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\] vssd1
+ vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\] vssd1
+ vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\] vssd1
+ vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net626 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout631 net633 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
X_09918_ _02829_ _02837_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout642 net644 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout653 net655 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08156__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 _04818_ vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__buf_2
XANTENNA__07307__S net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout675 net681 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__buf_2
Xfanout686 net687 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11337__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout697 net700 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
X_09849_ _04834_ _05520_ _05786_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07903__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ net1341 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09522__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09105__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11811_ _06637_ net456 net328 net1976 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791_ net1415 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11353__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14530_ clknet_leaf_130_wb_clk_i _02294_ _00895_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11742_ net2011 net266 net342 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__mux2_1
XANTENNA__11463__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15213__1578 vssd1 vssd1 vccd1 vccd1 _15213__1578/HI net1578 sky130_fd_sc_hd__conb_1
XANTENNA__08864__C1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11072__B net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14461_ clknet_leaf_60_wb_clk_i _02225_ _00826_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06875__D1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ net2212 net263 net349 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13412_ net1422 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input90_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ net1764 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] net836 vssd1 vssd1 vccd1
+ vccd1 _02504_ sky130_fd_sc_hd__mux2_1
X_14392_ clknet_leaf_8_wb_clk_i _02156_ _00757_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11499__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13343_ net1293 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ net1134 _06296_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08092__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13274_ net1401 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ net115 net1025 net902 net1731 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15013_ clknet_leaf_62_wb_clk_i _02733_ _01378_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__dfrtp_1
X_12225_ net1599 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09041__C1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09493__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net1712 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06910__A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ net829 _06523_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__and2_2
X_12087_ net615 _06653_ net457 net444 net1930 vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11247__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11038_ net1038 net831 net270 net668 vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11151__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09647__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ net1382 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11263__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14728_ clknet_leaf_15_wb_clk_i _02492_ _01093_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07122__A2 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14659_ clknet_leaf_25_wb_clk_i _02423_ _01024_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ _03140_ _03141_ net737 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\]
+ net948 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07131_ net750 _03072_ net1158 vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14382__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11202__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ net729 _03003_ _03002_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__o21a_1
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput212 net212 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_3_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput223 net223 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
Xoutput234 net234 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput245 net245 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput256 net256 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07594__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11438__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07964_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\]
+ net883 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09703_ net358 _05385_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a21o_1
XANTENNA__11157__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\] net793
+ net730 _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__o211a_1
X_07895_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\]
+ net880 _03836_ net1127 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09886__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09634_ net566 _05493_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand2_1
XANTENNA__10496__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07897__B1 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ net1205 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10996__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07005__A_N _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ net579 _05506_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12269__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11173__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__mux2_1
X_09496_ _05436_ _05437_ net578 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__mux2_1
XANTENNA__08846__C1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\]
+ net954 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout807_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14725__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08378_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11748__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07329_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\]
+ net890 vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09810__A1 _02923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07098__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ _06175_ _06176_ net282 vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__mux2_1
XANTENNA__07821__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ _04383_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] net671 vssd1
+ vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12010_ _06760_ net464 net365 net2327 vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__a22o_1
Xfanout1404 net1405 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1415 net1432 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1426 net1431 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 _06816_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 net462 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13961_ clknet_leaf_59_wb_clk_i _01725_ _00326_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout494 net495 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11782__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13563__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ net1427 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13892_ clknet_leaf_20_wb_clk_i _01656_ _00257_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12843_ net1253 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12774_ net1416 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XANTENNA__08837__C1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14513_ clknet_leaf_102_wb_clk_i _02277_ _00878_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_48_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ net594 _06479_ net465 _06808_ net1827 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12907__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14444_ clknet_leaf_7_wb_clk_i _02208_ _00809_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11656_ net2738 _06469_ net348 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06905__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\] net2879 net835
+ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__mux2_1
X_14375_ clknet_leaf_65_wb_clk_i _02139_ _00740_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11587_ _06453_ net2792 net452 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10947__B1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13326_ net1279 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ net147 net1029 net1020 net1829 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold909 team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\] vssd1
+ vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ net1247 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
X_10469_ _02765_ team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _06281_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__12642__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12208_ net1603 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08331__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ net1309 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11372__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ net1686 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__A _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07328__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07680_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\] net739
+ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09350_ _03989_ _05149_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08301_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\] net941
+ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ net607 _05145_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08232_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\]
+ net957 net916 vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07410__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13772__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14898__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10982__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\] net949
+ net915 vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__o21a_1
XANTENNA__10938__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07114_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\] net773
+ net747 _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07803__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\] net766
+ net727 _04035_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11867__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ net1123 _02984_ _02983_ net1156 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14128__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__B _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1032_A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12552__A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08359__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout492_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07031__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\] net1057
+ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ net1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\]
+ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07084__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout757_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07878_ net820 _03815_ _03819_ net719 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__o31a_1
XANTENNA__08531__A1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ net555 _05365_ net571 vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__o21a_1
X_06829_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] vssd1 vssd1 vccd1 vccd1
+ _02772_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout924_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10011__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _03529_ _04267_ net541 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12091__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ net566 _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _06627_ net2780 net393 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12490_ net1248 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ net2580 net397 _06760_ net503 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09876__B1_N net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08598__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ clknet_leaf_113_wb_clk_i _01924_ _00525_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\]
+ sky130_fd_sc_hd__dfrtp_1
X_11372_ net501 net622 _06738_ net406 net2221 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13111_ net1416 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XANTENNA__11777__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ _05968_ _05970_ _06127_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07270__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10944__A3 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ clknet_leaf_17_wb_clk_i _01855_ _00456_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13042_ net1403 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XANTENNA_input53_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ _03901_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11078__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1201 net1203 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
Xfanout1212 team_03_WB.instance_to_wrap.core.decoder.inst\[16\] vssd1 vssd1 vccd1
+ vccd1 net1212 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10185_ _03430_ _06025_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1223 net1229 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_4
XANTENNA__09193__D _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1234 net1239 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_4
Xfanout1245 team_03_WB.instance_to_wrap.core.decoder.inst\[8\] vssd1 vssd1 vccd1 vccd1
+ net1245 sky130_fd_sc_hd__buf_4
Xfanout1256 net1258 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_4
XANTENNA__11106__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1267 net1269 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_4
X_14993_ clknet_leaf_125_wb_clk_i net41 _01358_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1278 net1280 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_4
Xfanout280 _06409_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
Xfanout291 _05891_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_4
Xfanout1289 net1295 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_2
X_13944_ clknet_leaf_10_wb_clk_i _01708_ _00309_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08522__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07722__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ clknet_leaf_110_wb_clk_i _01639_ _00240_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12826_ net1371 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12757_ net1260 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11708_ _06750_ net390 net347 net2156 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12688_ net1416 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ clknet_leaf_32_wb_clk_i _02191_ _00792_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06931__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _06713_ net389 net354 net2685 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10157__A _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08589__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14358_ clknet_leaf_85_wb_clk_i _02122_ _00723_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10396__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold706 net142 vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\] vssd1
+ vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08684__S1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\] vssd1
+ vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ net1286 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XANTENNA__07261__A1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold739 team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\] vssd1
+ vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
X_14289_ clknet_leaf_94_wb_clk_i _02053_ _00654_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10148__A1 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14420__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ net1216 _04788_ _04789_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__nand3_1
XANTENNA__11896__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08761__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\] net774
+ net747 _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__o211a_1
X_08781_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\]
+ net974 net1071 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11138__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07732_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\] net789
+ _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14570__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08297__A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07663_ net1078 net885 team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\]
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09402_ _03641_ _05162_ net605 vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07594_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\]
+ net782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\] net749
+ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _05240_ _05274_ _05271_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__or3b_1
XFILLER_0_118_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08277__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _03682_ _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08215_ _04084_ _04155_ _04156_ _04154_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__o31a_1
XANTENNA__11170__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__B1 _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09195_ net548 _04825_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__nor2_1
XANTENNA__10067__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout505_A _06448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1247_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08146_ _02799_ _02801_ _02810_ _02812_ net1069 vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__a221o_4
XANTENNA__11584__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07788__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11597__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07252__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\]
+ net890 _04018_ net1119 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__o311a_1
XFILLER_0_60_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07028_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\]
+ net877 _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11336__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10006__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\] vssd1
+ vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14913__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08752__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\] vssd1
+ vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08752__B2 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 team_03_WB.instance_to_wrap.core.register_file.registers_state\[12\] vssd1
+ vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ net865 _04920_ _04915_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__o21ai_1
Xhold44 team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\] vssd1
+ vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\] vssd1
+ vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\] vssd1
+ vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\] vssd1
+ vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold88 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\] vssd1
+ vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ net272 net2807 net450 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__mux2_1
Xhold99 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\] vssd1
+ vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11345__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ net686 _05746_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ clknet_leaf_118_wb_clk_i _01424_ _00025_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10872_ net494 net594 _06469_ net521 net2147 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a32o_1
XANTENNA__11064__C net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12611_ net1296 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ net1282 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11361__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ net1385 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11080__B net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12473_ net1356 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15119__1500 vssd1 vssd1 vccd1 vccd1 _15119__1500/HI net1500 sky130_fd_sc_hd__conb_1
X_14212_ clknet_leaf_15_wb_clk_i _01976_ _00577_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11424_ _06517_ _06751_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nor2_1
X_15192_ net910 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14443__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07779__C1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14143_ clknet_leaf_114_wb_clk_i _01907_ _00508_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07243__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _06453_ net710 net695 vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] team_03_WB.instance_to_wrap.core.pc.current_pc\[22\]
+ _06146_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08991__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14074_ clknet_leaf_19_wb_clk_i _01838_ _00439_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11327__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286_ net513 net638 _06710_ net415 net2477 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a32o_1
XANTENNA_output257_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ net1265 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
X_10237_ _03602_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11878__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11239__C _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1021 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08743__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1031 _06283_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_2
Xfanout1042 net1043 vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_4
X_10168_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] net673 vssd1 vssd1 vccd1
+ vccd1 _06010_ sky130_fd_sc_hd__nand2_1
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__clkbuf_4
Xfanout1064 _02790_ vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07951__C1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11536__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__B _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1086 net1088 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__clkbuf_4
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_4
X_14976_ clknet_leaf_54_wb_clk_i _02728_ _01341_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dfrtp_1
X_10099_ _02832_ net314 _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__or3b_1
XFILLER_0_136_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11255__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ clknet_leaf_66_wb_clk_i _01691_ _00292_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07703__C1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10853__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06860__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13858_ clknet_leaf_132_wb_clk_i _01622_ _00223_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12809_ net1255 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12367__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ clknet_leaf_77_wb_clk_i _01553_ _00154_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11271__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11802__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09471__A2 _04149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07482__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ _03934_ _03941_ _03925_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10369__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11566__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold503 team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\] vssd1
+ vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold514 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\] vssd1
+ vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\] vssd1
+ vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\] vssd1
+ vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\] vssd1
+ vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11210__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14936__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _03169_ net662 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold558 team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\] vssd1
+ vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\] vssd1
+ vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08902_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\]
+ net959 net1067 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _05596_ _05633_ _05823_ _05611_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09082__S1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__A1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _02953_ net577 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nand2_4
Xhold1203 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\] vssd1
+ vssd1 vccd1 vccd1 net2787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\] vssd1
+ vssd1 vccd1 vccd1 net2798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\] vssd1
+ vssd1 vccd1 vccd1 net2809 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout288_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__C1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08739__B net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\] vssd1
+ vssd1 vccd1 vccd1 net2820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12041__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1247 team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\] vssd1
+ vssd1 vccd1 vccd1 net2831 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
Xhold1258 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\] vssd1
+ vssd1 vccd1 vccd1 net2842 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\] vssd1
+ vssd1 vccd1 vccd1 net2853 sky130_fd_sc_hd__dlygate4sd3_1
X_07715_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\]
+ net978 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\] net938
+ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout455_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07646_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\]
+ net788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\] net742
+ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10844__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07577_ net1128 _03515_ _03516_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout622_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__B _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11181__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09998__A0 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ net572 _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14466__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _03428_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ _05110_ _05113_ _05117_ _05119_ net558 net567 vssd1 vssd1 vccd1 vccd1 _05120_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout991_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08648__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__C net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08129_ _04069_ _04070_ net609 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_2
XANTENNA__07225__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08422__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08973__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ net1040 net833 net302 net666 vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__and4_1
XANTENNA__09864__A2_N _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11071_ _06613_ net2790 net421 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput101 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08725__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ net88 net87 vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14830_ clknet_leaf_61_wb_clk_i net1842 _01195_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ clknet_leaf_17_wb_clk_i _02525_ _01126_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11973_ net642 _06750_ net482 net372 net2076 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11790__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[9\] net314 net311 net321
+ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__and4_1
X_13712_ clknet_leaf_81_wb_clk_i _01476_ _00077_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14692_ clknet_leaf_42_wb_clk_i _02456_ _01057_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10835__A2 _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12037__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13643_ net1313 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_10855_ net827 _06453_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__and2_2
XFILLER_0_116_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10048__B1 _05907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11091__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13574_ net1424 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10786_ net314 net312 net323 vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__and3_1
XANTENNA__11522__C net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10599__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12525_ net1319 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11260__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12456_ net1340 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08604__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ net302 net2793 net401 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15175_ net1556 vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_2
XANTENNA__11012__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12387_ net1267 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
X_14126_ clknet_leaf_71_wb_clk_i _01890_ _00491_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11338_ net505 net629 _06721_ net406 net1826 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14057_ clknet_leaf_57_wb_clk_i _01821_ _00422_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\]
+ sky130_fd_sc_hd__dfrtp_1
X_15099__1480 vssd1 vssd1 vccd1 vccd1 _15099__1480/HI net1480 sky130_fd_sc_hd__conb_1
XANTENNA__09943__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11269_ net711 net271 net823 vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__and3_1
XANTENNA__08716__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ net1431 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10170__A _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ clknet_leaf_33_wb_clk_i _02711_ _01324_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10287__A0 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08480_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\] net942
+ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__o221a_1
XANTENNA__10826__A2 _06429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07431_ net1138 _03362_ _03372_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11205__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07362_ net1130 _03301_ _03302_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08101__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\] net954
+ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__or2_1
XANTENNA__07455__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07293_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__or3_1
XANTENNA__12825__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\]
+ net981 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08514__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 team_03_WB.instance_to_wrap.CPU_DAT_I\[9\] vssd1 vssd1 vccd1 vccd1 net1884
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 net177 vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold322 _02577_ vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold333 net199 vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08955__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 team_03_WB.instance_to_wrap.CPU_DAT_I\[13\] vssd1 vssd1 vccd1 vccd1 net1928
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08955__B2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\] vssd1
+ vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold366 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\] vssd1
+ vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold377 team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\] vssd1
+ vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 _02849_ vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_2
Xhold388 team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\] vssd1
+ vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _05871_ net1956 net294 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
Xhold399 team_03_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 net1983
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout813 _02847_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1112_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout824 _06558_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10999__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net849 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07654__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _03947_ net540 _04984_ _03944_ _02804_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__o32ai_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__buf_4
Xhold1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\] vssd1
+ vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net871 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_4
XANTENNA_hold1220_A team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout879 net882 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_4
Xhold1011 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\] vssd1
+ vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 team_03_WB.instance_to_wrap.ADR_I\[12\] vssd1 vssd1 vccd1 vccd1 net2606
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1033 team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\] vssd1
+ vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ net1216 _04755_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__or2_1
X_09796_ _05113_ _05130_ net558 vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__mux2_1
Xhold1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\] vssd1
+ vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1055 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\] vssd1
+ vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\] vssd1
+ vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\] vssd1
+ vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__a221o_1
Xhold1088 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\] vssd1
+ vssd1 vccd1 vccd1 net2672 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\] vssd1
+ vssd1 vccd1 vccd1 net2683 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09132__A1 _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__B2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__inv_2
XANTENNA__07143__B1 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ net1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\]
+ net872 net1144 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11115__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net1155 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] net842 vssd1 vssd1 vccd1
+ vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ net1953 net535 net596 _05881_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11242__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__D net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09840__C1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12310_ net1343 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07829__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ net1332 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09199__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ net1701 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09199__B2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08946__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net1707 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08946__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07267__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11950__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net2424 net419 _06636_ net507 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11054_ net510 net654 _06604_ net426 net1969 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07057__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11702__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _05890_ net1916 net288 vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14813_ clknet_leaf_61_wb_clk_i net1906 _01178_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14744_ clknet_leaf_117_wb_clk_i _02508_ _01109_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11956_ net627 _06733_ net466 net370 net2150 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a32o_1
XANTENNA__06908__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10907_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\] net313 net311 net322
+ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__and4_1
XANTENNA__07685__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14675_ clknet_leaf_54_wb_clk_i _02439_ _01040_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11887_ net619 _06696_ net458 net377 net2391 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a32o_1
XANTENNA__07685__B2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ net1310 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
X_10838_ net315 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__o31a_1
XFILLER_0_131_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11769__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07437__A1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13557_ net1430 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
X_10769_ net527 _06378_ _06379_ net532 net1896 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a32o_1
XFILLER_0_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12508_ net1341 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
X_13488_ net1334 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XANTENNA__08334__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14011__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12439_ net1414 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XANTENNA__10165__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15158_ net1539 vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13476__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ clknet_leaf_66_wb_clk_i _01873_ _00474_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\]
+ net900 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__or3_1
XFILLER_0_107_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15089_ net1470 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__09673__B _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06931_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\]
+ net773 net1123 vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__mux4_1
XANTENNA__07905__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09650_ _05356_ _05547_ _05589_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__o211a_1
XANTENNA__08796__S0 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ _02799_ _02801_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__nand2_8
XFILLER_0_101_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11427__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08601_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\] net996 net937
+ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__o221a_1
X_09581_ _05521_ _05522_ net577 vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ _04468_ _04473_ net870 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08463_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\] net914
+ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11472__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ net725 _03353_ _03354_ net1106 vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08394_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__o221a_1
XANTENNA__11162__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07345_ net1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\]
+ net885 vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1062_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07979__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07649__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\]
+ net777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\] net732
+ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o221a_1
X_09015_ _04895_ _04956_ net559 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1327_A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold130 team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\] vssd1
+ vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_83_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold141 team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\] vssd1
+ vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07087__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 team_03_WB.instance_to_wrap.ADR_I\[28\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\] vssd1
+ vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\] vssd1
+ vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07600__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\] vssd1
+ vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 team_03_WB.instance_to_wrap.CPU_DAT_I\[16\] vssd1 vssd1 vccd1 vccd1 net1780
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout610 net613 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
Xfanout621 net623 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09917_ _05082_ _05852_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__or3_1
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_2
Xfanout643 net644 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09889__C1 _05830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout954_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 _04818_ vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_4
Xfanout676 net681 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11337__C _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout687 net688 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_2
X_09848_ net540 _05787_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__o21a_1
XANTENNA__07364__B1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout698 net700 vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _04649_ _04956_ net563 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09105__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11810_ _06636_ net468 net329 net2434 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12790_ net1343 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A0 _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11353__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11741_ net1904 net267 net342 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__mux2_1
XANTENNA__07667__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11463__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__C net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06875__C1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ net2646 _06631_ net349 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
X_14460_ clknet_leaf_127_wb_clk_i _02224_ _00825_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13411_ net1421 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07419__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10623_ net1601 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\] net836 vssd1 vssd1 vccd1
+ vccd1 _02505_ sky130_fd_sc_hd__mux2_1
X_14391_ clknet_leaf_73_wb_clk_i _02155_ _00756_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13342_ net1292 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
X_10554_ team_03_WB.instance_to_wrap.BUSY_O team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ net604 net1137 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input83_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10974__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ net1396 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
X_10485_ net1989 net1025 net905 team_03_WB.instance_to_wrap.ADR_I\[21\] vssd1 vssd1
+ vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08919__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15012_ clknet_leaf_124_wb_clk_i net60 _01377_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12224_ net1750 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10726__A1 _05611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ net1724 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06910__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _06519_ net2517 net422 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
XANTENNA__07294__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12086_ net617 _06652_ net456 net444 net1931 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__a32o_1
XFILLER_0_60_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11037_ net2772 net426 _06594_ net507 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a22o_1
XANTENNA__11247__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07355__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11544__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08329__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__B1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09647__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__C1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ net1341 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
XANTENNA__12100__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14727_ clknet_leaf_118_wb_clk_i _02491_ _01092_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11454__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _06632_ net2638 net375 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__mux2_1
XANTENNA__07658__B2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__A _03136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ clknet_leaf_127_wb_clk_i _02422_ _01023_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_90_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ net1281 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
X_14589_ clknet_leaf_62_wb_clk_i _02353_ _00954_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07130_ net1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\]
+ net881 _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07469__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07061_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\] vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
XANTENNA__07830__A1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08999__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput213 net213 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
Xoutput224 net224 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput235 net235 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA__10717__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__B2 team_03_WB.instance_to_wrap.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput246 net246 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput257 net912 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XANTENNA__07594__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08791__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ net1099 net897 team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__o21a_1
XANTENNA__11438__B net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06914_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\]
+ net895 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09702_ _05073_ _05506_ _05638_ _04777_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\]
+ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__and2_1
XANTENNA__11157__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07897__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09633_ net585 _04775_ _05570_ _05573_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o311a_1
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06845_ net1200 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__inv_2
XANTENNA__11693__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout270_A _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _04269_ _04386_ _04448_ _04534_ net562 net565 vssd1 vssd1 vccd1 vccd1 _05506_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_78_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08239__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08515_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\]
+ net970 vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11173__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11445__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _05377_ _05381_ net567 vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__mux2_1
XANTENNA__08846__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout535_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1277_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08446_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\] net914
+ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o221a_1
XANTENNA__09859__A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08763__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078__1459 vssd1 vssd1 vccd1 vccd1 _15078__1459/HI net1459 sky130_fd_sc_hd__conb_1
X_08377_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\]
+ net961 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A _06559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07328_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\] net1119
+ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07379__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08074__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09810__A2 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\]
+ net774 net1124 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__mux4_1
XANTENNA__10009__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _05975_ _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11905__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1405 net1406 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__clkbuf_4
Xfanout1416 net1418 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1427 net1428 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _04075_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08003__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 _06816_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout462 net464 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ clknet_leaf_35_wb_clk_i _01724_ _00325_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_2
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11133__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 net498 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ net1388 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07888__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ clknet_leaf_24_wb_clk_i _01655_ _00256_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11684__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12842_ net1248 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12773_ net1271 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10644__A0 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08932__S0 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14512_ clknet_leaf_81_wb_clk_i _02276_ _00877_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\]
+ sky130_fd_sc_hd__dfrtp_1
X_11724_ net2041 net273 net341 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__A _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14443_ clknet_leaf_37_wb_clk_i _02207_ _00808_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\]
+ sky130_fd_sc_hd__dfrtp_1
X_11655_ net2777 _06454_ net348 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06905__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11303__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10606_ net2859 net2047 net835 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ net274 net2617 net453 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__mux2_1
X_14374_ clknet_leaf_79_wb_clk_i _02138_ _00739_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07499__S0 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10537_ net158 net1030 net1021 net1703 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13325_ net1318 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07812__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10468_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] _06280_ net680 vssd1
+ vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
X_13256_ net1342 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06921__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12207_ net1591 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__clkbuf_1
X_13187_ net1296 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
X_10399_ _06004_ _06069_ _06079_ _06078_ _03602_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o32a_1
XANTENNA__11372__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07228__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ net1607 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09009__A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12069_ _06631_ net2671 net363 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07328__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09443__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07752__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08300_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\] net925
+ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09280_ _05217_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08583__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08231_ net1058 _04171_ _04172_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13917__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08162_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\] net995
+ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07113_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\]
+ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\]
+ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__and2_1
XANTENNA__07803__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07044_ net1110 _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09556__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12044__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1025_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220__1580 vssd1 vssd1 vccd1 vccd1 _15220__1580/HI net1580 sky130_fd_sc_hd__conb_1
XANTENNA__11902__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _04935_ _04936_ net863 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__B _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08758__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07877_ net748 _03816_ _03818_ net804 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout652_A _06457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1394_A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ net561 _05357_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
XANTENNA__10874__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06828_ team_03_WB.instance_to_wrap.core.pc.current_pc\[24\] vssd1 vssd1 vccd1 vccd1
+ _02771_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ net566 _05486_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout917_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ net544 _04476_ _05101_ net561 vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08429_ _04369_ _04370_ net1210 vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11440_ net652 _06567_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09101__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11371_ net709 net298 net696 vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ _05968_ _05970_ _06127_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or3_1
XANTENNA__09528__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110_ net1343 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14090_ clknet_leaf_9_wb_clk_i _01854_ _00455_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13041_ net1315 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XANTENNA__11359__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ _04235_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] net670 vssd1
+ vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11354__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07558__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11078__B net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10184_ _03430_ _06025_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__and2_1
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input46_A gpio_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1213 net1217 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11793__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1235 net1236 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__clkbuf_4
Xfanout1246 team_03_WB.instance_to_wrap.core.decoder.inst\[7\] vssd1 vssd1 vccd1 vccd1
+ net1246 sky130_fd_sc_hd__buf_4
XANTENNA__09771__B _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14992_ clknet_leaf_124_wb_clk_i net40 _01357_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1257 net1258 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__buf_4
Xfanout270 _06509_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout1268 net1269 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_4
Xfanout1279 net1280 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__buf_4
Xfanout281 _06405_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 net295 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ clknet_leaf_86_wb_clk_i _01707_ _00308_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ clknet_leaf_100_wb_clk_i _01638_ _00239_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07730__B1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12825_ net1357 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ net1320 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12082__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11707_ _06749_ net389 net346 net1984 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ net1388 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08038__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14426_ clknet_leaf_7_wb_clk_i _02190_ _00791_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\]
+ sky130_fd_sc_hd__dfrtp_1
X_11638_ _06712_ net389 net354 net2467 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09786__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14357_ clknet_leaf_88_wb_clk_i _02121_ _00722_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ net508 net633 _06677_ net488 net1959 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold707 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\] vssd1
+ vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ net1284 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold718 team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\] vssd1
+ vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07747__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold729 team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\] vssd1
+ vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
X_14288_ clknet_leaf_113_wb_clk_i _02052_ _00653_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11269__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ net1418 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08746__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13484__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\]
+ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08780_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15077__1458 vssd1 vssd1 vccd1 vccd1 _15077__1458/HI net1458 sky130_fd_sc_hd__conb_1
XFILLER_0_100_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07731_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\] net763
+ net1037 vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09710__A1 _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11208__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09710__B2 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ net610 _03600_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11435__C net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ _05341_ _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07593_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\]
+ net782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\] net734
+ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11154__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15204__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ _05222_ _05236_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__or3b_1
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _03727_ _05147_ net606 vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09202__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08214_ net1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\]
+ net956 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\] net932
+ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08029__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09226__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09194_ net553 _04712_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11170__C net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ _02800_ _02802_ _02811_ _02813_ net1203 vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__o221a_2
XFILLER_0_31_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout400_A _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1142_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07788__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08076_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\]
+ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__or2_1
X_07027_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\]
+ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11336__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout867_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\] vssd1
+ vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\] vssd1
+ vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14395__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\] vssd1
+ vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _04916_ _04917_ _04919_ _04918_ net941 net861 vssd1 vssd1 vccd1 vccd1 _04920_
+ sky130_fd_sc_hd__mux4_1
Xhold45 team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\] vssd1
+ vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\] vssd1
+ vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_03_WB.instance_to_wrap.ADR_I\[24\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_93_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\] vssd1
+ vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ net743 _03867_ _03868_ _03869_ _03870_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__o32a_1
XANTENNA__11639__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\] vssd1
+ vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09162__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09701__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\] net308 net684 vssd1
+ vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__a21o_1
XANTENNA__11345__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07712__B1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ net827 _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__and2_2
XANTENNA__11064__D _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input100_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ net1348 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13590_ net1331 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11361__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11272__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ net1375 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11811__A2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09217__B1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12472_ net1368 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14211_ clknet_leaf_26_wb_clk_i _01975_ _00576_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11788__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ net297 net2758 net404 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15191_ net1572 vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_2
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14142_ clknet_leaf_49_wb_clk_i _01906_ _00507_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\]
+ sky130_fd_sc_hd__dfrtp_1
X_11354_ net502 net621 _06729_ net406 net2281 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07567__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10305_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] _06146_ vssd1 vssd1
+ vccd1 vccd1 _06147_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14073_ clknet_leaf_111_wb_clk_i _01837_ _00438_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\]
+ sky130_fd_sc_hd__dfrtp_1
X_11285_ net712 _06527_ net824 vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__and3_1
XANTENNA__14738__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10236_ _05068_ _02773_ net673 vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__mux2_1
X_13024_ net1407 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 _04085_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 net1022 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_4
X_10167_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__inv_2
Xfanout1032 net1033 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1043 _02791_ vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_8
Xfanout1054 _02791_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_4
Xfanout1065 net1068 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_4
Xfanout1076 _02789_ vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_4
X_14975_ clknet_leaf_31_wb_clk_i _02727_ _01340_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dfrtp_1
Xfanout1087 net1088 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13762__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10098_ _02924_ _02935_ _02936_ _05917_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a211o_1
Xfanout1098 net1105 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10838__B1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ clknet_leaf_79_wb_clk_i _01690_ _00291_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11255__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ clknet_leaf_4_wb_clk_i _01621_ _00222_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14118__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11552__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net1292 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13788_ clknet_leaf_119_wb_clk_i _01552_ _00153_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15211__1577 vssd1 vssd1 vccd1 vccd1 _15211__1577/HI net1577 sky130_fd_sc_hd__conb_1
XANTENNA__07467__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12739_ net1296 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09759__A1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13479__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ clknet_leaf_59_wb_clk_i _02173_ _00774_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07219__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11566__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08967__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold504 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\] vssd1
+ vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold515 team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\] vssd1
+ vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07865__S0 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold526 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\] vssd1
+ vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\] vssd1
+ vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\] vssd1
+ vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _05879_ net2245 net292 vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
Xhold559 team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\] vssd1
+ vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\]
+ net959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\] net1202
+ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__o221a_1
XFILLER_0_110_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09881_ _05803_ _05811_ _05821_ _05646_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__or4b_1
XANTENNA__08195__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08832_ net560 _04713_ _04773_ net574 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__o211a_1
Xhold1204 team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\] vssd1
+ vssd1 vccd1 vccd1 net2788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1215 team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\] vssd1
+ vssd1 vccd1 vccd1 net2799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_03_WB.instance_to_wrap.ADR_I\[31\] vssd1 vssd1 vccd1 vccd1 net2810
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\] vssd1
+ vssd1 vccd1 vccd1 net2821 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ net1214 _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or2_1
Xhold1248 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\] vssd1
+ vssd1 vccd1 vccd1 net2832 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1259 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1 net2843
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07714_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\] net789
+ net1011 _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08694_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\]
+ net978 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\] net922
+ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07645_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\]
+ net788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\] vssd1
+ vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1092_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07576_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\]
+ net897 _03517_ net1147 vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__o311a_1
XFILLER_0_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11181__B net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ net607 _05124_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__nor2_1
XANTENNA__11254__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10078__A _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout615_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1357_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09246_ _03391_ _05152_ net605 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09586__B _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ net547 net357 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11401__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08128_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] net1017 net682 vssd1
+ vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08958__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07818__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08059_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\]
+ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11070_ net827 net279 vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11059__D net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput102 wbs_we_i vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_10021_ net84 net83 net86 net85 vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__or4_1
XANTENNA__10532__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07933__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14760_ clknet_leaf_118_wb_clk_i _02524_ _01125_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09686__B1 _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ net636 _06749_ net477 net371 net2389 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a32o_1
XANTENNA__07850__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13711_ clknet_leaf_98_wb_clk_i _01475_ _00076_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10923_ net315 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[9\]
+ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__o31a_1
X_14691_ clknet_leaf_42_wb_clk_i _02455_ _01056_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ net1309 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ _06450_ _06451_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_71_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11091__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14410__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ net1402 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11522__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10785_ _06381_ _06382_ _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__or3b_2
XFILLER_0_32_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12524_ net1304 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08661__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15076__1457 vssd1 vssd1 vccd1 vccd1 _15076__1457/HI net1457 sky130_fd_sc_hd__conb_1
XFILLER_0_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12455_ net1389 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10716__A _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11548__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ _06434_ net2733 net404 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__mux2_1
XANTENNA__08413__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15174_ net1555 vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_2
XFILLER_0_133_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ net1353 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14125_ clknet_leaf_110_wb_clk_i _01889_ _00490_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\]
+ sky130_fd_sc_hd__dfrtp_1
X_11337_ net1242 net832 _06413_ net666 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14056_ clknet_leaf_34_wb_clk_i _01820_ _00421_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ net518 net641 _06701_ net415 net2538 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ net1410 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10219_ _06024_ _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nor2_1
X_11199_ net281 net2605 net492 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10523__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__B1 _03865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09017__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14958_ clknet_leaf_56_wb_clk_i _02710_ _01323_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09677__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07760__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07688__C1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ clknet_leaf_87_wb_clk_i _01673_ _00274_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\]
+ sky130_fd_sc_hd__dfrtp_1
X_14889_ clknet_leaf_44_wb_clk_i _02652_ _01254_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12378__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07430_ net1130 _03367_ _03369_ _03371_ net720 vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__o41a_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12028__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11236__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07361_ net816 _03290_ net717 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08101__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09100_ net440 net431 _05041_ net554 vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07292_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\]
+ net777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\] net1126
+ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08591__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09031_ _04971_ _04972_ net862 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__o21a_1
XANTENNA__10087__B_N _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__B2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__A1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold301 _02580_ vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07838__S0 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 team_03_WB.instance_to_wrap.ADR_I\[0\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold323 team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\] vssd1
+ vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07000__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold334 team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\] vssd1
+ vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__C1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold345 _02584_ vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold356 net200 vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold367 team_03_WB.instance_to_wrap.CPU_DAT_I\[24\] vssd1 vssd1 vccd1 vccd1 net1951
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold378 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\] vssd1
+ vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 team_03_WB.instance_to_wrap.core.ru.state\[6\] vssd1 vssd1 vccd1 vccd1 net1973
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _03821_ net661 vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout803 net805 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout825 net826 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10999__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout398_A _06757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__clkbuf_4
X_09864_ _03947_ _04984_ _05805_ _02945_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12052__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout847 net849 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__buf_8
Xfanout858 _04083_ vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_4
XANTENNA__10514__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07915__B1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_8
Xhold1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\] vssd1
+ vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11711__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1105_A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\] vssd1
+ vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08815_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\] net1060
+ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a221o_1
Xhold1023 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\] vssd1
+ vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ net579 _05736_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or2_1
Xhold1034 team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\] vssd1
+ vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout565_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\] vssd1
+ vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07391__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1056 team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\] vssd1
+ vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1067 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\] vssd1
+ vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__a221o_1
Xhold1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\] vssd1
+ vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\] vssd1
+ vssd1 vccd1 vccd1 net2673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07670__A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09132__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ _04607_ _04618_ net848 vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__mux2_8
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12288__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11192__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__or3_1
XANTENNA__07694__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11227__A0 _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07559_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\] vssd1
+ vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10570_ net1783 net538 net599 _05880_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08643__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08643__B2 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_750 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09229_ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__inv_2
XANTENNA__07851__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12240_ net1839 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08006__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12171_ net1752 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11950__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11122_ net281 net653 net705 net699 vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold890 team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\] vssd1
+ vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11367__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ net1040 net833 _06536_ net669 vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__and4_2
XFILLER_0_21_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07057__S1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07906__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ _05889_ net1886 net288 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07283__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__C1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14812_ clknet_leaf_41_wb_clk_i net1677 _01177_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07580__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ clknet_leaf_11_wb_clk_i _02507_ _01108_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11955_ net616 _06732_ net457 net369 net2182 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a32o_1
XANTENNA__06908__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ net315 _05846_ net320 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14674_ clknet_leaf_54_wb_clk_i _02438_ _01039_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11886_ net622 _06695_ net462 net378 net1819 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__a32o_1
XANTENNA__14926__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11218__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13625_ net1421 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10837_ net302 net2556 net521 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__mux2_1
XANTENNA__12926__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13556_ net1429 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ _05142_ net603 vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09831__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12507_ net1364 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07842__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ net1397 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10699_ _05455_ _06310_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12438_ net1343 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15157_ net1538 vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
X_12369_ net1303 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14108_ clknet_leaf_119_wb_clk_i _01872_ _00473_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07070__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15088_ net1469 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11277__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ net1147 net1159 vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__or2_4
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14039_ clknet_leaf_86_wb_clk_i _01803_ _00404_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09898__B1 _05403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14456__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08796__S1 _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ _02800_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__nor2_2
XANTENNA__07373__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13492__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\]
+ net973 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XANTENNA__07912__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09580_ _05396_ _05402_ net567 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08531_ net1213 _04471_ _04472_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11457__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08322__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11216__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ net931 _04402_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11209__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07413_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\] net738
+ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__o221a_1
X_08393_ net1238 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\]
+ net991 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\] net1074
+ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07344_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\] net724
+ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09210__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07275_ net1132 _03216_ net722 vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12047__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout313_A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1055_A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09014_ _04923_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08389__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold120 _02573_ vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09050__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold131 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[13\] vssd1 vssd1 vccd1
+ vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\] vssd1
+ vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 _02631_ vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\] vssd1
+ vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\] vssd1
+ vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 net141 vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold197 _02587_ vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 _06295_ vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_2
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
X_09916_ _02837_ _05142_ _05799_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__or4b_1
XFILLER_0_22_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout622 net626 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
Xfanout633 net645 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout655 _06457_ vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
XANTENNA__09880__A _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout666 _06564_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_4
Xfanout677 net681 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
XANTENNA__11696__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ net572 _04739_ net665 _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
Xfanout688 net689 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_2
XANTENNA__11337__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15075__1456 vssd1 vssd1 vccd1 vccd1 _15075__1456/HI net1456 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _05270_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08729_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07116__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11740_ net594 net263 net469 _06808_ net1893 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a32o_1
XANTENNA__08864__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11353__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11671_ net2110 net264 net349 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ net1400 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08077__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10622_ net1729 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] net837 vssd1 vssd1 vccd1
+ vccd1 _02506_ sky130_fd_sc_hd__mux2_1
XANTENNA__08435__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08616__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14390_ clknet_leaf_85_wb_clk_i _02154_ _00755_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10959__C1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11620__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ net1286 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ team_03_WB.instance_to_wrap.core.ru.state\[0\] team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nor2_1
XANTENNA__07824__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08092__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14329__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10974__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input76_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ net1401 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
X_10484_ net1900 net1027 net904 team_03_WB.instance_to_wrap.ADR_I\[22\] vssd1 vssd1
+ vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11796__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ clknet_leaf_126_wb_clk_i net59 _01376_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13577__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ net1680 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09041__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A0 _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07575__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12154_ net1714 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08170__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11097__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _06628_ net2137 net422 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12085_ net619 _06651_ net458 net444 net1799 vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11687__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ net631 _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__nor2_1
XANTENNA__11151__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ net1344 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08304__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14726_ clknet_leaf_123_wb_clk_i _02490_ _01091_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11938_ net263 net2615 net376 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ clknet_leaf_134_wb_clk_i _02421_ _01022_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11869_ net269 net2065 net382 vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__mux2_1
XANTENNA__06961__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ net1327 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08068__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14588_ clknet_leaf_126_wb_clk_i _02352_ _00953_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_32_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13539_ net1271 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11611__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07060_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\]
+ net796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\] net743
+ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__a221o_1
XANTENNA__09965__A _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07291__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13487__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15209_ net910 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput214 net214 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput225 net225 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
Xoutput236 net236 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_50_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput247 net247 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput258 net258 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__08240__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07594__A1 net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11390__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07962_ net610 _03900_ _03902_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08218__S0 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13846__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__C net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ _02954_ _04477_ _05126_ _05640_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a311o_1
X_06913_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\] net773
+ net747 _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__o211a_1
XANTENNA__11678__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\]
+ net880 _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11142__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] _02803_ net539 _05571_
+ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__o2bb2a_1
X_06844_ net1185 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09205__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09099__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _05178_ _05180_ _05503_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
XANTENNA__11173__C net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ net574 _05383_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
XANTENNA__08846__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10653__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11850__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\] net931
+ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout430_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09859__B _05746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1172_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\]
+ net961 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
XANTENNA__08255__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11602__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07327_ _03265_ _03268_ net816 vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09810__A3 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07258_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\] net1148
+ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o221a_1
XANTENNA__07821__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout897_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09023__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\]
+ net754 vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
XANTENNA__11905__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__A2 _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1406 net1433 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__buf_2
Xfanout1417 net1418 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1428 net1431 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__buf_4
XFILLER_0_100_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout430 net436 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08003__B _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout452 _06801_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 net464 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07337__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 net485 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11133__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout485 _06800_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ net1336 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
Xfanout496 net498 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13890_ clknet_leaf_130_wb_clk_i _01654_ _00255_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14001__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ net1247 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10892__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[15\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12094__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12772_ net1314 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XANTENNA__08298__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14511_ clknet_leaf_97_wb_clk_i _02275_ _00876_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ net594 _06469_ net459 _06808_ net2035 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11841__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08932__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__B _05106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ clknet_leaf_2_wb_clk_i _02206_ _00807_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\]
+ sky130_fd_sc_hd__dfrtp_1
X_11654_ net2357 _06620_ net352 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10605_ net1971 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] net836 vssd1 vssd1 vccd1
+ vccd1 _02523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14373_ clknet_leaf_107_wb_clk_i _02137_ _00738_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07499__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ net301 net2853 net453 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10947__A2 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ net1283 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10536_ net161 net1030 net1021 net1909 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13255_ net1403 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10724__A _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _02775_ _06279_ net285 vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13869__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ net1593 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08222__C1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13186_ net1348 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
X_10398_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] _06141_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07576__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11372__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ net1665 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10580__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ net264 net2661 net363 vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__mux2_1
XANTENNA__07328__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ net1243 net828 _06478_ net667 vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12085__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10635__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14709_ clknet_leaf_118_wb_clk_i _02473_ _01074_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\]
+ net955 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\] net932
+ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14644__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08161_ _04095_ _04102_ net867 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07112_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\] net793
+ net730 _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08092_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\] net764
+ net740 _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a211o_1
XANTENNA__11060__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15074__1455 vssd1 vssd1 vccd1 vccd1 _15074__1455/HI net1455 sky130_fd_sc_hd__conb_1
XANTENNA__08461__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07043_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\]
+ net773 net1123 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13010__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07016__B1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09556__A2 _05485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11899__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ net1209 _04932_ _04933_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__nand3_1
XANTENNA__10571__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_A _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\] net788 net743
+ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout380_A _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__C _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout478_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\] net780
+ net729 _03817_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09615_ _04778_ _05551_ _05555_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_1294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11184__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06827_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] vssd1 vssd1 vccd1 vccd1
+ _02770_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1387_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12076__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net570 _05487_ net326 vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08819__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11823__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout812_A _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _05415_ _05418_ net566 vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11404__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12091__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\] net934
+ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08359_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\] net935
+ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07255__B1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ net502 net623 _06737_ net405 net2240 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06151_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\]
+ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07270__A3 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13040_ net1429 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__inv_2
XANTENNA__11359__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08014__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07102__S0 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ _04619_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] net672 vssd1
+ vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1203 net1207 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
XANTENNA__10562__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
XANTENNA__08949__A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1225 net1228 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09544__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1236 net1238 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__buf_2
Xfanout1247 net1251 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_4
XANTENNA_input39_A gpio_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ clknet_leaf_6_wb_clk_i net39 _01356_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout1258 net1270 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_2
Xfanout271 _06491_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_2
Xfanout1269 net1270 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
XANTENNA__11375__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13942_ clknet_leaf_93_wb_clk_i _01706_ _00307_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09180__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ clknet_leaf_96_wb_clk_i _01637_ _00238_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07621__A1_N net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12067__A0 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ net1368 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_104_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__A2_N _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10617__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12755_ net1259 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10719__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11706_ _06748_ net388 net347 net1840 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ net1341 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14425_ clknet_leaf_111_wb_clk_i _02189_ _00790_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\]
+ sky130_fd_sc_hd__dfrtp_1
X_11637_ _06711_ net388 net355 net2577 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a22o_1
XANTENNA__08669__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11042__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14356_ clknet_leaf_91_wb_clk_i _02120_ _00721_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11568_ net2368 net488 _06797_ net511 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ net1284 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
Xhold708 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\] vssd1
+ vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire683 _02933_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_1
X_10519_ net148 net1023 net1019 net1797 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
Xhold719 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\] vssd1
+ vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ clknet_leaf_99_wb_clk_i _02051_ _00652_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ _06620_ net2764 net394 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13238_ net1338 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XANTENNA__11269__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11984__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13169_ net1315 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XANTENNA__11896__A3 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11285__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _03670_ _03671_ net1154 vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09710__A2 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ net610 _03601_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07182__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11435__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09400_ _03352_ _04475_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12058__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ _03531_ _03533_ net810 vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10608__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09331_ _05230_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09262_ _05198_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11820__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08213_ net1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\]
+ net955 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\] net916
+ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09226__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09193_ net548 net441 net433 _04739_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__or4_1
XFILLER_0_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10067__C net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__B1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _02799_ _02801_ _02810_ _02812_ net1043 vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a221o_2
XANTENNA__08533__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07788__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08985__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12055__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ _04010_ _04011_ _04016_ net1153 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1135_A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\]
+ net877 _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout595_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11336__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1302_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold13 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\] vssd1
+ vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_03_WB.instance_to_wrap.ADR_I\[10\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout762_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\] vssd1
+ vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\] vssd1
+ vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\] vssd1
+ vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\]
+ net893 net1121 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a211o_1
Xhold68 _02627_ vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold79 team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\] vssd1
+ vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07859_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _06465_ _06466_ _06467_ net586 vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__o211a_4
X_15189__1570 vssd1 vssd1 vccd1 vccd1 _15189__1570/HI net1570 sky130_fd_sc_hd__conb_1
XFILLER_0_116_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09529_ _05469_ _05470_ net565 vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11272__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ net1350 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XANTENNA__08673__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08009__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ net1414 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XANTENNA__12754__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ clknet_leaf_127_wb_clk_i _01974_ _00575_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ net270 net2597 net401 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__mux2_1
X_15190_ net1571 vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07779__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14141_ clknet_leaf_66_wb_clk_i _01905_ _00506_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[495\]
+ sky130_fd_sc_hd__dfrtp_1
X_11353_ net274 net709 net696 vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10783__B1 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07059__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] team_03_WB.instance_to_wrap.core.pc.current_pc\[20\]
+ _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and3_1
X_14072_ clknet_leaf_118_wb_clk_i _01836_ _00437_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11284_ net517 net642 _06709_ net416 net2376 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13023_ net1375 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
X_10235_ _06073_ _06074_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10535__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11878__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1000 net1001 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1011 _02869_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_8
Xfanout1022 _06286_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
X_10166_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or2_1
Xfanout1033 net1034 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07951__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1044 net1045 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1055 net1057 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_4
XANTENNA__11309__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1066 net1068 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
Xfanout1077 _02788_ vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_8
XFILLER_0_22_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14974_ clknet_leaf_62_wb_clk_i _02726_ _01339_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dfrtp_1
Xfanout1088 _02787_ vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_4
X_10097_ _02832_ _02926_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_117_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ clknet_leaf_109_wb_clk_i _01689_ _00290_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15073__1454 vssd1 vssd1 vccd1 vccd1 _15073__1454/HI net1454 sky130_fd_sc_hd__conb_1
XANTENNA__07703__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08900__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13856_ clknet_leaf_133_wb_clk_i _01620_ _00221_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06927__A net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ net1399 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09303__A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13787_ clknet_leaf_26_wb_clk_i _01551_ _00152_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\]
+ sky130_fd_sc_hd__dfrtp_1
X_10999_ net1039 net832 net278 net668 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__and4_2
XFILLER_0_123_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11271__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12738_ net1348 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
XANTENNA__10168__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11979__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12669_ net1381 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
XANTENNA__12664__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14408_ clknet_leaf_27_wb_clk_i _02172_ _00773_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09759__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08967__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ clknet_leaf_18_wb_clk_i _02103_ _00704_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold505 team_03_WB.instance_to_wrap.ADR_I\[14\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\] vssd1
+ vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07865__S1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06978__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold527 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\] vssd1
+ vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold538 team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\] vssd1
+ vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold549 net191 vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08900_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\]
+ net959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\] net1067
+ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__o221a_1
XANTENNA__13495__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__inv_2
XANTENNA__10526__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08831_ net564 _04740_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or3_1
Xhold1205 team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\] vssd1
+ vssd1 vccd1 vccd1 net2789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07942__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1216 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\] vssd1
+ vssd1 vccd1 vccd1 net2800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11219__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\] vssd1
+ vssd1 vccd1 vccd1 net2811 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__mux2_1
Xhold1238 team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\] vssd1
+ vssd1 vccd1 vccd1 net2822 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1249 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\] vssd1
+ vssd1 vccd1 vccd1 net2833 sky130_fd_sc_hd__dlygate4sd3_1
X_07713_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__or3_1
XANTENNA__10829__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ net940 _04633_ _04634_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07644_ net812 _03577_ net720 vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\]
+ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1085_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _04711_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07458__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11254__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09245_ _05185_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12574__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09176_ net439 net431 _05041_ net547 vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08958__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ net721 _04041_ _04047_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o31a_2
XFILLER_0_86_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10094__A _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08058_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout977_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ net1018 _02943_ _02947_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10517__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08499__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08186__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ net74 net77 net76 net75 vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__or4b_2
XFILLER_0_60_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07933__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11971_ net632 _06748_ net469 net372 net2236 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a32o_1
XANTENNA__09686__B2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ clknet_leaf_70_wb_clk_i _01474_ _00075_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10922_ net686 _05706_ _06401_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__a21oi_1
X_14690_ clknet_leaf_53_wb_clk_i _02454_ _01055_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10835__A4 _06403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13641_ net1396 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09679__A1_N _05568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10853_ net691 _05623_ net586 vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12037__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__A0 _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10048__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13572_ net1329 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XANTENNA__08646__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10784_ _06393_ _06391_ _06392_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__and3b_4
XANTENNA__08110__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11799__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12523_ net1257 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07578__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ net1411 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11548__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11405_ net276 net2648 net404 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15173_ net1554 vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_2
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12385_ net1291 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14124_ clknet_leaf_4_wb_clk_i _01888_ _00489_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11336_ net504 net624 _06720_ net406 net2382 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a32o_1
XFILLER_0_120_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ clknet_leaf_66_wb_clk_i _01819_ _00420_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11267_ net1243 net834 net300 net669 vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__and4_2
XANTENNA__10508__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07517__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09374__B1 _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ net1339 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
X_10218_ _06057_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__and2_1
XANTENNA__11547__B _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] _06394_ _06455_ vssd1
+ vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nand3_4
XANTENNA__07924__A1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ _03138_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14957_ clknet_leaf_61_wb_clk_i _02709_ _01322_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07137__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11563__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ clknet_leaf_92_wb_clk_i _01672_ _00273_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07688__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__C1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14888_ clknet_leaf_44_wb_clk_i _02651_ _01253_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13839_ clknet_leaf_97_wb_clk_i _01603_ _00204_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11236__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07360_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08101__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07291_ _03229_ _03232_ net819 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10907__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[12\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11502__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10995__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\]
+ net981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\] net944
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07488__A team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07860__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11539__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__C1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 net210 vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07838__S1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold313 team_03_WB.instance_to_wrap.ADR_I\[16\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold324 team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\] vssd1
+ vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_03_WB.instance_to_wrap.CPU_DAT_I\[14\] vssd1 vssd1 vccd1 vccd1 net1919
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\] vssd1
+ vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\] vssd1
+ vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _05870_ net1800 net292 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
Xhold368 _02595_ vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold379 team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\] vssd1
+ vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_2
XANTENNA__08168__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout815 _02847_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout826 _06558_ vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__buf_4
XANTENNA__09208__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10999__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__clkbuf_4
X_09863_ _03947_ _04984_ net541 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o21a_1
XANTENNA__08112__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net849 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 _04083_ vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__clkbuf_8
X_08814_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\]
+ net976 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__mux2_1
Xhold1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\] vssd1
+ vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\] vssd1
+ vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ _05084_ _05091_ _05117_ _05086_ net562 net570 vssd1 vssd1 vccd1 vccd1 _05736_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1000_A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\] vssd1
+ vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1035 team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\] vssd1
+ vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\] vssd1
+ vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1057 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\] vssd1
+ vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net860 _04685_ _04686_ _04684_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1068 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\] vssd1
+ vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10788__S net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout460_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07128__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\] vssd1
+ vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09668__B2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08258__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _04610_ _04611_ _04617_ _04614_ net1060 net1077 vssd1 vssd1 vccd1 vccd1 _04618_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08340__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__B2 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ net1166 net872 team_03_WB.instance_to_wrap.core.register_file.registers_state\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__a21o_1
XANTENNA__11192__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12019__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout725_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _03496_ _03499_ net819 vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08782__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09840__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07489_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11412__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _04532_ _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07851__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14878__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ net437 net429 _04503_ net550 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__o31a_1
XFILLER_0_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15072__1453 vssd1 vssd1 vccd1 vccd1 _15072__1453/HI net1453 sky130_fd_sc_hd__conb_1
XFILLER_0_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12170_ net1726 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08721__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11121_ _06449_ net627 _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__or3_4
XANTENNA__14108__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\] vssd1
+ vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold891 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\] vssd1
+ vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ net508 net655 _06603_ net427 net1860 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a32o_1
XANTENNA__08022__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__C1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ _05888_ net1730 net287 vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__mux2_1
XANTENNA__11702__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ clknet_leaf_60_wb_clk_i net1872 _01176_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11383__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ net615 _06731_ net457 net369 net2480 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a32o_1
X_14742_ clknet_leaf_116_wb_clk_i _02506_ _01107_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10905_ net691 _05697_ net586 vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__o21a_1
X_14673_ clknet_leaf_55_wb_clk_i _02437_ _01038_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net624 _06694_ net463 net377 net2287 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13624_ net1316 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10836_ _06436_ _06437_ _06435_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11769__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13555_ net1329 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
XANTENNA__08095__B1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10767_ team_03_WB.instance_to_wrap.core.pc.current_pc\[0\] net603 vssd1 vssd1 vccd1
+ vccd1 _06378_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09292__C1 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__C_N net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11322__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13103__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12506_ net1365 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07842__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13486_ net1392 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ net1736 net531 net526 _06336_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ net1268 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10729__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15156_ net1537 vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ net1428 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ clknet_leaf_30_wb_clk_i _01871_ _00472_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\]
+ sky130_fd_sc_hd__dfrtp_1
X_11319_ _06626_ net2735 net409 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07070__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15087_ net1468 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
X_12299_ net1253 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168__1549 vssd1 vssd1 vccd1 vccd1 _15168__1549/HI net1549 sky130_fd_sc_hd__conb_1
X_14038_ clknet_leaf_93_wb_clk_i _01802_ _00403_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09898__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07358__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 _02802_ sky130_fd_sc_hd__nand3b_2
XANTENNA__08867__A _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08570__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__A2 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ net1059 _04469_ _04470_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__or3_1
XANTENNA__11457__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08858__C1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08461_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\] net952 net914
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07412_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\]
+ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08392_ net861 _04330_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07343_ net738 _03281_ _03282_ _03283_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__o32a_1
XFILLER_0_50_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09822__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09210__B _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07274_ _02872_ _03214_ _03215_ _02870_ _03213_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08107__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09013_ net443 net435 _04953_ net547 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07011__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08389__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07946__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\] vssd1
+ vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 net208 vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold132 team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\] vssd1
+ vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06850__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold143 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[26\] vssd1 vssd1 vccd1
+ vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold154 team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\] vssd1
+ vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11468__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\] vssd1
+ vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12063__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\] vssd1
+ vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07600__A3 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1215_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 _02585_ vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _06295_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\] vssd1
+ vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 net613 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_4
X_09915_ _05646_ _05676_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__and3_1
Xfanout623 net626 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_2
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07349__C1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout645 _06458_ vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_4
Xfanout656 net658 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_4
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout667 _06564_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_4
XANTENNA__08010__B1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ net543 _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand2_1
Xfanout678 net680 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08561__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 _02840_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09777_ _05240_ _05241_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11407__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08728_ net1213 _04668_ _04669_ _04665_ _04667_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09510__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08659_ net860 _04599_ _04600_ _04598_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11670_ net2543 _06630_ net351 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ net2353 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] net837 vssd1 vssd1 vccd1
+ vccd1 _02507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09813__B2 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ net1284 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
X_10552_ net1136 _06293_ _06292_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07824__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13271_ net1401 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10974__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10483_ net118 net1026 net902 net1787 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_129_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15010_ clknet_leaf_41_wb_clk_i net58 _01375_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12222_ net1685 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input69_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11384__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ net1776 vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07052__B2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11104_ net829 net297 vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__and2_2
XANTENNA__11097__B net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ net623 _06650_ net461 net447 net1854 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14080__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11035_ net716 _06503_ net701 vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__or3_1
XANTENNA__13648__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11317__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11439__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__S1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ net1373 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08304__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ clknet_leaf_123_wb_clk_i _02489_ _01090_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_11937_ _06631_ net2811 net375 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__mux2_1
XANTENNA__11263__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14656_ clknet_leaf_134_wb_clk_i _02420_ _01021_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11868_ _06527_ net2187 net382 vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06961__S1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09311__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ net314 net312 net323 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__a31o_1
X_13607_ net1280 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XANTENNA__08068__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_24 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14587_ clknet_leaf_32_wb_clk_i _02351_ _00952_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\]
+ sky130_fd_sc_hd__dfstp_1
X_11799_ net2523 _06628_ net334 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07815__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13538_ net1279 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10176__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11987__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13469_ net1394 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
XANTENNA__09965__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07830__A3 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15208_ net1576 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_112_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput215 net215 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput226 net226 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput237 net237 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10192__A _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ net1520 vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
Xoutput248 net248 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput259 net259 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_107_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08791__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07961_ net610 _03900_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__a21o_1
XANTENNA__08791__B2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08218__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11438__D net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ _03866_ _05012_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06912_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\]
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07892_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[335\]
+ net1149 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21o_1
XANTENNA__14573__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _03314_ _04415_ net663 _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06843_ net1156 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__clkinv_4
XANTENNA__07897__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13008__A net1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _05180_ _05503_ _05178_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__o21ai_1
X_08513_ net870 _04451_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__or3_1
X_15071__1452 vssd1 vssd1 vccd1 vccd1 _15071__1452/HI net1452 sky130_fd_sc_hd__conb_1
X_09493_ net582 _05433_ _05434_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11173__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08444_ net544 _04384_ _04355_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06845__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12058__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout423_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07326_ net801 _03266_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07806__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07379__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10086__B _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09008__C1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07257_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\]
+ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1332_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07676__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07188_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\]
+ net755 vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
XANTENNA__11366__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1407 net1409 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__buf_4
Xfanout1418 net1432 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__buf_2
Xfanout420 _06635_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_4
Xfanout431 net432 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1429 net1430 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11669__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout453 _06801_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout464 net485 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07337__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 net477 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__clkbuf_4
Xfanout486 _06779_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_2
X_09829_ _05263_ _05264_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07888__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12840_ net1293 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10892__A2 _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12771_ net1302 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14510_ clknet_leaf_68_wb_clk_i _02274_ _00875_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\]
+ sky130_fd_sc_hd__dfrtp_1
X_11722_ _06454_ net594 net458 _06808_ net1834 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09131__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14441_ clknet_leaf_57_wb_clk_i _02205_ _00806_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\]
+ sky130_fd_sc_hd__dfrtp_1
X_15167__1548 vssd1 vssd1 vccd1 vccd1 _15167__1548/HI net1548 sky130_fd_sc_hd__conb_1
XFILLER_0_83_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11653_ net2284 _06619_ net348 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09798__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ net1836 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] net836 vssd1 vssd1 vccd1
+ vccd1 _02524_ sky130_fd_sc_hd__mux2_1
X_14372_ clknet_leaf_20_wb_clk_i _02136_ _00737_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ net302 net2532 net452 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13323_ net1288 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
X_10535_ net162 net1029 net1020 net1871 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11600__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13254_ net1429 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
X_10466_ _06047_ _06049_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__xnor2_1
X_12205_ net1659 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13185_ net1258 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
XANTENNA__08222__B1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10397_ _06222_ _06223_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] net677
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12136_ net1719 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11109__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12067_ _06630_ net2702 net364 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11018_ net494 net646 _06582_ net425 net2012 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09306__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08210__A net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12085__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_max_cap590_A _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ net1251 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14708_ clknet_leaf_120_wb_clk_i _02472_ _01073_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14639_ clknet_leaf_98_wb_clk_i _02403_ _01004_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_56_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08160_ net1208 _04100_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07111_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08091_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\]
+ net875 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__and3_1
XANTENNA__11060__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11510__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07042_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\] vssd1
+ vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11348__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07016__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08213__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11899__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08993_ net1055 _04934_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10571__B2 _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15218__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07944_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__D _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07875_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\]
+ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout373_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06826_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] vssd1 vssd1 vccd1 vccd1
+ _02769_ sky130_fd_sc_hd__inv_2
X_09614_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] _02803_ net540 _05553_
+ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10874__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _05413_ _05417_ net562 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10796__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout540_A _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09476_ _05416_ _05417_ net556 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11823__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07170__S net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\]
+ net965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\] net918
+ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout805_A _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\] net917
+ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__o221a_1
XANTENNA__11587__A0 _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07309_ net1109 _03249_ _03250_ net1119 vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13201__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] net675 _06157_ _06160_
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _06091_ _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12000__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11359__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10011__A0 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08755__A1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] _02819_ _06023_ vssd1
+ vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10562__B2 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1216 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
Xfanout1226 net1228 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__clkbuf_4
Xfanout1237 net1238 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14990_ clknet_leaf_124_wb_clk_i net38 _01355_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1248 net1250 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_4
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
Xfanout272 _06483_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
XANTENNA__11375__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout283 net286 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
X_13941_ clknet_leaf_87_wb_clk_i _01705_ _00306_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_4
X_13872_ clknet_leaf_82_wb_clk_i _01636_ _00237_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12823_ net1417 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XANTENNA__11391__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ net1420 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
XANTENNA__09483__A2 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ _06747_ net389 net346 net1958 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ net1319 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14424_ clknet_leaf_2_wb_clk_i _02188_ _00789_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\]
+ sky130_fd_sc_hd__dfrtp_1
X_11636_ _06710_ net391 net354 net2463 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11578__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A3 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08669__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11042__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14355_ clknet_leaf_110_wb_clk_i _02119_ _00720_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11567_ net637 net706 net268 net697 vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11330__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ net149 net1023 net1019 net1858 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__a22o_1
X_13306_ net1292 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14286_ clknet_leaf_70_wb_clk_i _02050_ _00651_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\] vssd1
+ vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ _06619_ net2417 net393 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__mux2_1
XANTENNA__07747__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13986__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13237_ net1263 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
X_10449_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] _06265_ net679 vssd1
+ vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
X_15070__1451 vssd1 vssd1 vccd1 vccd1 _15070__1451/HI net1451 sky130_fd_sc_hd__conb_1
XANTENNA__11269__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__A0 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08746__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13168_ net1429 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
XANTENNA__11750__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net238 net99 net101 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__and3b_1
X_13099_ net1257 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XANTENNA__11285__B _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07660_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07182__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07591_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\] net782
+ net733 _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12397__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09330_ _04646_ _05229_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11805__A1 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09261_ _05201_ _05202_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08212_ _04152_ _04153_ net856 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09192_ _05130_ _05133_ net557 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08814__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11569__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__D net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07237__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _02800_ _02802_ _02811_ _02813_ net1223 vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__o221a_2
XFILLER_0_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08074_ net740 _04012_ _04013_ _04014_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o32a_1
X_07025_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\]
+ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08737__A1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08198__C1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09645__S net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\] vssd1
+ vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08976_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\]
+ net985 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__mux2_1
X_15166__1547 vssd1 vssd1 vccd1 vccd1 _15166__1547/HI net1547 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 _02613_ vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold36 team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\] vssd1
+ vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\] vssd1
+ vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ net1089 net893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\]
+ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o21a_1
Xhold58 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\] vssd1
+ vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\] vssd1
+ vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07858_ net1149 _03798_ _03799_ net820 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__o31a_1
XFILLER_0_98_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07789_ _03729_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06920__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11415__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__S0 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09528_ _05348_ _05352_ net561 vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07476__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ net548 _04712_ _05132_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08673__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11361__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ net1348 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
XANTENNA__08724__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07228__A1 _03169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ net2444 net403 _06754_ net508 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10232__B1 _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14140_ clknet_leaf_120_wb_clk_i _01904_ _00505_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11352_ net504 net624 _06728_ net405 net1949 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07567__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11980__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10783__A1 _02842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] team_03_WB.instance_to_wrap.core.pc.current_pc\[18\]
+ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14071_ clknet_leaf_86_wb_clk_i _01835_ _00436_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ net713 net296 net825 vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__and3_1
XANTENNA__08728__A1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ net1378 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
X_10234_ _06073_ _06074_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__nor2_1
XANTENNA_input51_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07936__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1001 net1010 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_2
XFILLER_0_24_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1012 _02821_ vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__buf_4
X_10165_ _03724_ _06005_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1023 _06283_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_4
Xfanout1034 _05905_ vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__clkbuf_4
Xfanout1045 net1050 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_4
X_14973_ clknet_leaf_61_wb_clk_i _02725_ _01338_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dfrtp_1
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__buf_4
X_10096_ net314 _05429_ _05936_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__or4_1
XANTENNA__14634__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1078 net1088 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
Xfanout1089 net1092 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13924_ clknet_leaf_16_wb_clk_i _01688_ _00289_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08900__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ clknet_leaf_122_wb_clk_i _01619_ _00220_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06927__B net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13106__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ net1411 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14784__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ net2808 net427 _06571_ net518 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XANTENNA__09456__A2 _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13786_ clknet_leaf_8_wb_clk_i _01550_ _00151_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08113__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07467__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12737_ net1290 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ net1347 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XANTENNA__09957__C net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14407_ clknet_leaf_64_wb_clk_i _02171_ _00772_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07219__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _06693_ net388 net355 net2657 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XANTENNA__09759__A3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ net1415 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XANTENNA__08967__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11566__A3 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14338_ clknet_leaf_131_wb_clk_i _02102_ _00703_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold506 net213 vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 net216 vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 net224 vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold539 team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\] vssd1
+ vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14269_ clknet_leaf_68_wb_clk_i _02033_ _00634_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12680__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__S1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11723__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ net442 net434 _04770_ _03105_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o31a_1
XFILLER_0_42_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1206 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\] vssd1
+ vssd1 vccd1 vccd1 net2790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\] vssd1
+ vssd1 vccd1 vccd1 net2801 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\] net1060
+ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__a221o_1
Xhold1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\] vssd1
+ vssd1 vccd1 vccd1 net2812 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\] vssd1
+ vssd1 vccd1 vccd1 net2823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11446__D net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09144__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07712_ _03652_ _03653_ net1154 vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__o21a_1
XANTENNA__10829__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\] net977 net922
+ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__a221o_1
XANTENNA__07155__B1 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07643_ net816 _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__nand2_1
XANTENNA__11743__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A1_N net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07574_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\]
+ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09313_ net580 _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07458__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08655__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11254__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_A _06810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09244_ _04119_ _05184_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1078_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _05115_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12066__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08126_ net1139 _04057_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08958__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09080__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10765__A1 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11962__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07630__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ _03995_ _03998_ net817 vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1412_A net1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07008_ _02949_ _02947_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08959_ net852 _04899_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or3_1
X_11970_ net637 _06747_ net478 net371 net2341 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__A2 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08343__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ net270 net2367 net521 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__mux2_1
XANTENNA__07850__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13640_ net1315 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
X_10852_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[20\] net308 net684 vssd1
+ vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14037__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13571_ net1308 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XANTENNA__08646__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10783_ _02842_ _05918_ _06385_ _06293_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08110__A2 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07859__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ net1257 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input99_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12453_ net1288 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XANTENNA__14187__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11404_ net278 net2672 net402 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ net1553 vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_2
XANTENNA__09071__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12384_ net1408 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08413__A3 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11953__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14123_ clknet_leaf_18_wb_clk_i _01887_ _00488_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\]
+ sky130_fd_sc_hd__dfrtp_1
X_11335_ _06409_ net710 net695 vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ net515 net634 _06700_ net416 net2258 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a32o_1
X_14054_ clknet_leaf_81_wb_clk_i _01818_ _00419_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11705__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ _06024_ _06058_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nor2_1
X_13005_ net1301 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ net2261 net420 _06679_ net517 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__a22o_1
XANTENNA__07385__B1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__A2 _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10148_ _04207_ net670 _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09126__A1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14956_ clknet_leaf_63_wb_clk_i _02708_ _01321_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10079_ _05921_ _05922_ net316 _05920_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__a211o_1
XANTENNA__07137__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__A2 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ clknet_leaf_110_wb_clk_i _01671_ _00272_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11563__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07688__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14887_ clknet_leaf_43_wb_clk_i _02650_ _01252_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13838_ clknet_leaf_71_wb_clk_i _01602_ _00203_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10894__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ clknet_leaf_67_wb_clk_i _01533_ _00134_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10444__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07290_ net803 _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__or3_1
XANTENNA__10995__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15165__1546 vssd1 vssd1 vccd1 vccd1 _15165__1546/HI net1546 sky130_fd_sc_hd__conb_1
XANTENNA__08591__C _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10747__A1 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11944__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\] vssd1
+ vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold314 _02619_ vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 team_03_WB.instance_to_wrap.CPU_DAT_I\[3\] vssd1 vssd1 vccd1 vccd1 net1909
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09600__A_N _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold336 team_03_WB.instance_to_wrap.ADR_I\[6\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\] vssd1
+ vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold358 team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\] vssd1
+ vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 team_03_WB.instance_to_wrap.CPU_DAT_I\[17\] vssd1 vssd1 vccd1 vccd1 net1953
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _03312_ net660 vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout805 _02849_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout816 _02846_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_6
X_09862_ _05278_ _05281_ _05300_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__nand3_1
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_4
Xfanout838 _06304_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_4
Xfanout849 _04096_ vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07376__B1 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__B2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\]
+ net976 vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__mux2_1
XANTENNA__07009__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\] vssd1
+ vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\] vssd1
+ vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _05421_ _05734_ net576 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__mux2_2
Xhold1025 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\] vssd1
+ vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1036 team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\] vssd1
+ vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\] vssd1
+ vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\] vssd1
+ vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\] net923
+ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07128__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\] vssd1
+ vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06848__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07679__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08675_ _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout453_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1195_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10683__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07626_ net1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__or3_1
XANTENNA__11192__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07557_ net803 _03497_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08628__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout620_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net821 vssd1 vssd1 vccd1
+ vccd1 _03430_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09227_ _03280_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07851__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09158_ net570 _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10738__A1 _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__A0 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08109_ net727 _04048_ _04049_ net1108 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__a31o_1
XANTENNA__07603__A1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09089_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\] net918
+ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08800__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11120_ net1038 net700 vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11950__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\] vssd1
+ vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\] vssd1
+ vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold892 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\] vssd1
+ vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ net705 net269 net826 vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__and3_2
XANTENNA__11367__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _05887_ net1832 net289 vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__mux2_1
XANTENNA__07906__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07462__S0 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ clknet_leaf_56_wb_clk_i net1910 _01175_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08316__C1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09134__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ clknet_leaf_117_wb_clk_i _02505_ _01106_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11383__B _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07580__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ net619 _06730_ net458 net369 net2000 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10904_ net299 net2159 net524 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__mux2_1
X_14672_ clknet_leaf_52_wb_clk_i _02436_ _01037_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ net630 _06693_ net468 net380 net2224 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13623_ net1404 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10835_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[23\] _05865_ net321 _06403_
+ net687 vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11603__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13554_ net1421 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ net2080 net532 net527 _06377_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09831__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ net1354 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
XANTENNA__07842__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ _06317_ _06333_ _06335_ net604 vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__o2bb2a_1
X_13485_ net1392 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12436_ net1321 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XANTENNA__11926__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07055__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ net1536 vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12367_ net1407 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ clknet_leaf_23_wb_clk_i _01870_ _00471_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07528__S net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ _06625_ net2829 net410 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09309__A _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15086_ net1467 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
X_12298_ net1256 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11249_ net275 net713 net825 vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__and3_1
X_14037_ clknet_leaf_87_wb_clk_i _01801_ _00402_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11277__C _06509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10889__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__A1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12103__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11293__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14939_ clknet_leaf_40_wb_clk_i _02694_ _01304_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11457__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08460_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XANTENNA__14352__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07411_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or3_1
X_08391_ net852 _04331_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__or3_1
XANTENNA__09807__C1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11513__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07342_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\]
+ net885 net1115 vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08086__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11090__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\]
+ net777 vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 net173 vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[16\] vssd1
+ vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold122 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\] vssd1
+ vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 team_03_WB.instance_to_wrap.ADR_I\[2\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold155 team_03_WB.instance_to_wrap.core.ru.state\[2\] vssd1 vssd1 vccd1 vccd1 net1739
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\] vssd1
+ vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 net165 vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\] vssd1
+ vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 team_03_WB.instance_to_wrap.CPU_DAT_I\[18\] vssd1 vssd1 vccd1 vccd1 net1783
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 net603 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_2
X_09914_ _05659_ _05822_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout613 _02842_ vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1110_A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07349__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout624 net626 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__C _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__B2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout635 net645 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1208_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08546__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout646 net648 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_4
XANTENNA__08010__A1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_2
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ net573 _04739_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__or2_1
XANTENNA__11696__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout570_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _06563_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__buf_4
Xfanout679 net680 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_2
XANTENNA__11484__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07364__A3 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _05709_ _05712_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__or3_4
XFILLER_0_20_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06988_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] _02827_ _02829_ vssd1
+ vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\] net937
+ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__A0 team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\] net924
+ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07609_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\]
+ net782 vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__mux2_1
XANTENNA__06875__A2 team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08589_ net863 _04530_ _04525_ net846 vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__o211a_1
XANTENNA__10828__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11423__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08077__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10620_ net2844 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] net836 vssd1 vssd1 vccd1
+ vccd1 _02508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09813__A2 _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ net1135 _06293_ _06292_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07824__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11620__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09828__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14995__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ net119 net1027 net904 net1651 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
X_13270_ net1338 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ net1765 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07037__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11384__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08785__C1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net1721 vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08033__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _06627_ net2687 net421 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12083_ _06787_ net467 net444 net1892 vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08537__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11034_ net2246 net425 _06592_ net501 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XANTENNA__08001__A1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11687__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15164__1545 vssd1 vssd1 vccd1 vccd1 _15164__1545/HI net1545 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11439__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12985_ net1356 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10647__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ clknet_leaf_15_wb_clk_i _02488_ _01089_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12100__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09799__A _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ net264 net2787 net375 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14655_ clknet_leaf_109_wb_clk_i _02419_ _01020_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11867_ net296 net2302 net383 vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13606_ net1280 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08068__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ net692 _05541_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14586_ clknet_leaf_21_wb_clk_i _02350_ _00951_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\]
+ sky130_fd_sc_hd__dfstp_1
X_11798_ net2569 _06627_ net336 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09804__A2 _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07276__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13537_ net1283 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10749_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] net602 vssd1 vssd1 vccd1
+ vccd1 _06367_ sky130_fd_sc_hd__or2_1
XANTENNA__11611__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15000__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13468_ net1393 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XANTENNA__06951__A team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08642__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15207_ net910 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09568__B2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ net1300 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_13399_ net1395 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
XANTENNA__07579__B1 _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput216 net216 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput227 net227 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XANTENNA__08776__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput238 net238 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
X_15138_ net1519 vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XANTENNA__08240__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput249 net249 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15069_ net1450 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
X_07960_ net613 _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08528__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09473__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ net1147 net883 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nand2_1
X_07891_ net803 _03828_ _03831_ _03832_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__a22o_1
XANTENNA__11678__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11508__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net541 _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nand2_1
XANTENNA__10886__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09740__A1 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06842_ net1148 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__clkinv_4
XANTENNA__08089__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ _05308_ _05501_ _05182_ _05190_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10638__A0 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ _04452_ _04453_ net859 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09492_ _05313_ _05432_ _05320_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07503__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08443_ net545 _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13024__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08374_ net1199 _04312_ _04315_ net845 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__o31a_1
XANTENNA__08118__A net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07325_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\] net740
+ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1060_A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout416_A _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__C _05746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1158_A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10810__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07187_ net1106 _03123_ _03124_ _03126_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__o32a_1
XFILLER_0_108_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1325_A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11366__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1408 net1409 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__buf_4
Xfanout410 _06717_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1419 net1420 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__buf_4
XFILLER_0_100_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout421 net424 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout432 net436 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _04075_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout454 net455 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout465 net467 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10877__A0 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout476 net477 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ _05442_ _05669_ net578 vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__mux2_1
Xfanout487 _06779_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
Xfanout498 net505 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09759_ _03243_ net540 _04922_ _05700_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08917__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12770_ net1353 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XANTENNA__08298__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11721_ net2060 _06446_ net341 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11841__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14440_ clknet_leaf_34_wb_clk_i _02204_ _00805_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\]
+ sky130_fd_sc_hd__dfrtp_1
X_11652_ net2731 _06618_ net351 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08028__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ net1727 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] net838 vssd1 vssd1 vccd1
+ vccd1 _02525_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07258__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ clknet_leaf_24_wb_clk_i _02135_ _00736_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12773__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ net275 net2724 net455 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10801__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input81_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13322_ net1279 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ net163 net1024 net1022 net1676 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11389__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ net2871 net680 _06275_ _06278_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__o22a_1
X_13253_ net1271 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12204_ net1626 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08222__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10396_ net283 _06143_ _06220_ net677 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ net1409 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
X_12135_ net1625 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07576__A3 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08773__A2 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__B1 _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13765__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _06528_ net2813 net363 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11328__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11017_ net703 net273 net822 vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__and3_1
XANTENNA__10868__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07733__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12948__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12085__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ net1340 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
XANTENNA__08637__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ clknet_leaf_120_wb_clk_i _02471_ _01072_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09322__A _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _06620_ net2833 net374 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12899_ net1302 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14638_ clknet_leaf_68_wb_clk_i _02402_ _01003_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14569_ clknet_leaf_60_wb_clk_i _02333_ _00934_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07110_ _03050_ _03051_ net809 vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08090_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08461__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08461__B2 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10915__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07041_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\] net1148
+ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a221o_1
XANTENNA__11299__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11348__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14540__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08213__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08992_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\]
+ net954 net1069 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__mux4_1
XANTENNA__10931__A _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10571__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07943_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\] net743
+ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A1 _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07874_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\]
+ net780 vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09613_ _03280_ _04532_ net664 _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__a22o_1
X_06825_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] vssd1 vssd1 vccd1 vccd1
+ _02768_ sky130_fd_sc_hd__inv_2
XANTENNA__11184__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_A _06817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ _05405_ _05414_ net561 vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__mux2_1
XANTENNA__12076__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09232__A _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ net546 _04179_ _05083_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12069__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1275_A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ _04362_ _04367_ net868 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ net936 _04297_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07308_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\]
+ net765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\] net1154
+ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08282__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163__1544 vssd1 vssd1 vccd1 vccd1 _15163__1544/HI net1544 sky130_fd_sc_hd__conb_1
X_08288_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[887\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07239_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\] net1125
+ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__o221a_1
XFILLER_0_21_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10250_ _03426_ _06090_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13788__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10181_ _04646_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] net672 vssd1
+ vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10562__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1207 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_6
Xfanout1216 net1217 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_4
Xfanout1227 net1228 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_2
Xfanout1238 net1239 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09704__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout273 _06473_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__buf_2
X_13940_ clknet_leaf_92_wb_clk_i _01704_ _00305_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11375__C net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
Xfanout295 _05859_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09180__A2 _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ clknet_leaf_97_wb_clk_i _01635_ _00236_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07810__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12822_ net1343 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14413__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12753_ net1312 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11704_ _06746_ net389 net346 net2008 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
X_12684_ net1302 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ clknet_leaf_74_wb_clk_i _02187_ _00788_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11635_ _06709_ net391 net354 net2169 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07597__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ clknet_leaf_105_wb_clk_i _02118_ _00719_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08192__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ net506 net631 _06675_ net488 net2235 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13305_ net1284 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
X_10517_ net150 net1024 net1022 net1806 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
XANTENNA__07651__C1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14285_ clknet_leaf_104_wb_clk_i _02049_ _00650_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ _06618_ net2694 net394 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_113_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13236_ net1324 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10448_ _06264_ _06263_ net284 vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07403__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net1388 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
X_10379_ net283 _06207_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15052__1584 vssd1 vssd1 vccd1 vccd1 net1584 _15052__1584/LO sky130_fd_sc_hd__conb_1
X_12118_ net1136 net911 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__or2_1
XANTENNA__09317__A _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ net1248 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ _06618_ net2814 net364 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__mux2_1
XANTENNA__11285__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07182__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07590_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\]
+ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08367__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _05012_ _05200_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__nand2_1
XANTENNA__14906__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08891__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11018__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ net1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\] net955 net916
+ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09191_ _05131_ _05132_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ net1212 _02820_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nand2_4
XANTENNA__09631__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07300__A team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\]
+ net890 net1118 vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07024_ net746 _02964_ _02965_ net1156 vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a31o_1
XANTENNA__09926__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1023_A _06283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A1 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09227__A _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold15 team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\] vssd1
+ vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\] vssd1
+ vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[19\] vssd1 vssd1 vccd1
+ vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\]
+ net878 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold48 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[30\] vssd1 vssd1 vccd1
+ vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold59 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\] vssd1
+ vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__B1 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07970__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07857_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\]
+ net781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\] net1159
+ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout650_A _06457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout748_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__B1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10600__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07788_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\] net1122
+ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09527_ _05349_ _05360_ net555 vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__mux2_1
XANTENNA__08348__S1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08122__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09458_ _05129_ _05131_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _05306_ _05307_ _05311_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11431__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _06503_ _06751_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nor2_1
XANTENNA__13212__A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08425__A1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11351_ net301 net711 net696 vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__and3_1
XANTENNA__07633__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] team_03_WB.instance_to_wrap.core.pc.current_pc\[16\]
+ _06142_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__and3_1
X_14070_ clknet_leaf_84_wb_clk_i _01834_ _00435_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11282_ net512 net639 _06708_ net415 net1907 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13021_ net1366 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10233_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__inv_2
XANTENNA__10535__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07936__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11732__A1 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10164_ _03724_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input44_A gpio_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 net1010 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09137__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1024 _06283_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_2
Xfanout1035 net1036 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__clkbuf_4
Xfanout1046 net1047 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
X_14972_ clknet_leaf_56_wb_clk_i _02724_ _01337_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dfrtp_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10095_ _05435_ _05453_ _05518_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__or4b_1
XFILLER_0_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__clkbuf_4
Xfanout1079 net1088 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_2
XANTENNA__09153__A2 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13923_ clknet_leaf_18_wb_clk_i _01687_ _00288_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11606__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ clknet_leaf_78_wb_clk_i _01618_ _00219_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11248__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ net1275 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13785_ clknet_leaf_83_wb_clk_i _01549_ _00150_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08113__B1 net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ net641 _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__nor2_1
XANTENNA__09456__A3 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12736_ net1408 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XANTENNA__08664__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13953__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07872__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ net1360 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ clknet_leaf_77_wb_clk_i _02170_ _00771_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13122__A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08416__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ _06692_ net390 net355 net2465 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a22o_1
XANTENNA__09613__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ net1346 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14337_ clknet_leaf_2_wb_clk_i _02101_ _00702_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11549_ net498 net619 _06659_ net486 net1879 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a32o_1
XANTENNA__06978__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold507 team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\] vssd1
+ vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11971__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold518 team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\] vssd1
+ vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\] vssd1
+ vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14268_ clknet_leaf_128_wb_clk_i _02032_ _00633_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13219_ net1263 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14199_ clknet_leaf_87_wb_clk_i _01963_ _00564_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10526__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11723__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__A_N _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1207 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\] vssd1
+ vssd1 vccd1 vccd1 net2791 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ net1200 _04701_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2_1
Xhold1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\] vssd1
+ vssd1 vccd1 vccd1 net2802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\] vssd1
+ vssd1 vccd1 vccd1 net2813 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\] net1143
+ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10829__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\]
+ net978 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__mux2_1
X_15162__1543 vssd1 vssd1 vccd1 vccd1 _15162__1543/HI net1543 sky130_fd_sc_hd__conb_1
XFILLER_0_135_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07155__A1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11516__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07642_ net1107 _03582_ _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07573_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__or3_1
XANTENNA__09213__C net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ _02938_ _05125_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08655__A1 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ _04119_ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout329_A net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09174_ net439 net431 _05068_ net554 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__o31a_1
XFILLER_0_12_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11411__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08125_ net1133 _04062_ _04064_ _04066_ net721 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__o41a_1
XFILLER_0_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09080__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1140_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1238_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08056_ net801 _03996_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout698_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07007_ net1018 _02943_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1405_A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11714__A1 _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\] net941
+ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07909_ net732 _03849_ _03850_ net1112 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07146__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ net585 _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__nor2_1
XANTENNA__08343__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__A3 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _06507_ _06508_ _06506_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[20\] net306 vssd1
+ vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__nand2_1
XANTENNA__13976__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ net1313 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08646__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10782_ _06381_ _06382_ _06388_ net1136 vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ net1252 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
X_15051__1583 vssd1 vssd1 vccd1 vccd1 net1583 _15051__1583/LO sky130_fd_sc_hd__conb_1
XFILLER_0_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ net1298 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XANTENNA__07578__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11402__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ net303 net2732 net404 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
X_15171_ net1552 vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ net1354 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11953__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07875__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ clknet_leaf_3_wb_clk_i _01886_ _00487_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\]
+ sky130_fd_sc_hd__dfrtp_1
X_11334_ net507 net630 _06719_ net407 net2125 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14601__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ clknet_leaf_109_wb_clk_i _01817_ _00418_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ net716 net272 net826 vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__and3_1
XANTENNA__10508__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07909__B1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net1297 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
X_15109__1490 vssd1 vssd1 vccd1 vccd1 _15109__1490/HI net1490 sky130_fd_sc_hd__conb_1
X_10216_ _06023_ _03206_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11196_ net656 net707 net266 net698 vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10147_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] net670 vssd1 vssd1 vccd1
+ vccd1 _05989_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_48 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14751__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14955_ clknet_leaf_63_wb_clk_i _02707_ _01320_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07137__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _02937_ _05342_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13906_ clknet_leaf_103_wb_clk_i _01670_ _00271_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_14886_ clknet_leaf_51_wb_clk_i _02649_ _01251_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11563__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13837_ clknet_leaf_106_wb_clk_i _01601_ _00202_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ clknet_leaf_26_wb_clk_i _01532_ _00133_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09330__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ net1389 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XANTENNA__11641__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13699_ clknet_leaf_26_wb_clk_i _01463_ _00064_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11071__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10995__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__C net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07860__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09062__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11944__A1 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\] vssd1
+ vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 team_03_WB.instance_to_wrap.core.i_hit vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07612__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 _02574_ vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14281__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold337 _02609_ vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 team_03_WB.instance_to_wrap.ADR_I\[4\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09930_ _05869_ net2001 net292 vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold359 team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\] vssd1
+ vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08248__S0 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13849__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout806 net811 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_8
Xfanout817 _02846_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
X_09861_ _05802_ _05686_ _05676_ _05659_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_68_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout828 _06387_ vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
XANTENNA__07376__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08112__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
X_08812_ net869 _04753_ net847 vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a21oi_1
X_09792_ _05526_ _05600_ net570 vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__mux2_1
Xhold1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\] vssd1
+ vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\] vssd1
+ vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1026 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\] vssd1
+ vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1037 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\] vssd1
+ vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\] net939
+ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a221o_1
Xhold1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\] vssd1
+ vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\] vssd1
+ vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07128__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10132__A0 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\] net925
+ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07025__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07625_ _03529_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__nand2_1
XANTENNA__11880__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1090_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1188_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\]
+ net779 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\] net748
+ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09240__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__B2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__C1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ _03391_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout613_A _02842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1355_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _03314_ _05160_ net605 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10199__A0 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ _05095_ _05098_ net555 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08487__S0 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08108_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\] net740
+ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ _05028_ _05029_ net1210 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09534__B1_N _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\] net788
+ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold860 team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\] vssd1
+ vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\] vssd1
+ vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold882 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\] vssd1
+ vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap590 _02989_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__buf_4
XFILLER_0_25_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08013__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\] vssd1
+ vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ net2812 net426 _06602_ net513 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a22o_1
XANTENNA__11699__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__A1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _05886_ net2090 net287 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__mux2_1
XANTENNA__08022__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07462__S1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__A2 _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ clknet_leaf_120_wb_clk_i _02504_ _01105_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ net622 _06729_ net462 net370 net2553 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a32o_1
XANTENNA__11383__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11871__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10903_ net686 _06493_ _06494_ _06492_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__o31a_4
XFILLER_0_135_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14671_ clknet_leaf_55_wb_clk_i _02435_ _01036_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11883_ net640 _06692_ net481 net379 net2179 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14154__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13622_ net1422 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ net315 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[23\]
+ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__o31a_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09816__B1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13553_ net1429 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XANTENNA__11623__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10765_ team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] _05082_ net602 vssd1
+ vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__mux2_1
XANTENNA__09292__A1 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12504_ net1362 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
X_13484_ net1397 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10696_ _06312_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_129_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12435_ net1265 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15161__1542 vssd1 vssd1 vccd1 vccd1 _15161__1542/HI net1542 sky130_fd_sc_hd__conb_1
XANTENNA__10729__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07055__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15154_ net1535 vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ net1337 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
XANTENNA__08252__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14105_ clknet_leaf_103_wb_clk_i _01869_ _00470_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\]
+ sky130_fd_sc_hd__dfrtp_1
X_11317_ _06624_ net2782 net410 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15085_ net1466 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
X_12297_ net1252 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
X_14036_ clknet_leaf_92_wb_clk_i _01800_ _00401_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\]
+ sky130_fd_sc_hd__dfrtp_1
X_11248_ net519 net643 _06691_ net415 net2053 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a32o_1
XANTENNA__07358__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07358__B2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ net639 _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12103__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09044__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08858__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14938_ clknet_leaf_126_wb_clk_i _02693_ _01303_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11293__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11862__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14869_ clknet_leaf_53_wb_clk_i net1846 _01234_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07410_ _02782_ _03351_ net610 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__mux2_1
X_08390_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\] net942
+ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__o221a_1
XANTENNA__08375__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__A1 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ net1078 net885 team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\]
+ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10968__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07272_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\]
+ net779 vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ net844 _04931_ _04937_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a31o_4
XFILLER_0_54_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14797__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07046__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\] vssd1
+ vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08243__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\] vssd1
+ vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold123 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\] vssd1
+ vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\] vssd1
+ vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08794__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold145 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[7\] vssd1 vssd1 vccd1
+ vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[18\] vssd1 vssd1 vccd1
+ vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\] vssd1
+ vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 _02578_ vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09934__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _05854_ _05718_ _05697_ _05686_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__and4b_1
Xhold189 net219 vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 _06295_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_2
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__buf_2
XANTENNA__11145__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_A _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 net639 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
Xfanout647 net648 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_2
X_09844_ net583 _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nand2_1
X_15050__1582 vssd1 vssd1 vccd1 vccd1 net1582 _15050__1582/LO sky130_fd_sc_hd__conb_1
Xfanout658 _06457_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1103_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08641__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _06563_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_4
XANTENNA__09235__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ net358 _05485_ _05714_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout563_A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06987_ _02838_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\] net920
+ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11853__A0 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\] net940
+ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout730_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout828_A _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\]
+ net782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\] net734
+ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__o221a_1
XANTENNA__08285__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ _04526_ _04527_ _04529_ _04528_ net934 net858 vssd1 vssd1 vccd1 vccd1 _04530_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11605__A0 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10828__B _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07539_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\]
+ net795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\] net1148
+ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a221oi_1
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11005__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ team_03_WB.instance_to_wrap.core.d_hit net689 vssd1 vssd1 vccd1 vccd1 _06293_
+ sky130_fd_sc_hd__nor2_4
XFILLER_0_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09209_ _04073_ _05147_ net606 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_1
X_10481_ net120 net1027 net904 net2345 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ net1641 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07037__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11384__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12151_ net1672 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ net827 net270 vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ _06786_ net468 net445 net2155 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a22o_1
Xhold690 team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\] vssd1
+ vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08537__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net622 _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__nor2_1
XANTENNA__08001__A2 _02821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12097__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12984_ net1373 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11844__A0 _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14723_ clknet_leaf_123_wb_clk_i _02487_ _01088_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11935_ _06630_ net2506 net376 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09799__B _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14654_ clknet_leaf_57_wb_clk_i _02418_ _01019_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\]
+ sky130_fd_sc_hd__dfstp_1
X_11866_ _06683_ net476 net382 net1835 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a22o_1
X_13605_ net1282 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10817_ net303 net2658 net523 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14585_ clknet_leaf_111_wb_clk_i _02349_ _00950_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11797_ net2557 _06505_ net333 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07276__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13536_ net1280 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10748_ net2070 net532 net526 _06366_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13467_ net1393 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10679_ net604 _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06951__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ net912 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09568__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ net1374 vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13398_ net1308 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07766__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput217 net217 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XANTENNA__08776__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15137_ net1518 vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
Xoutput228 net228 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12349_ net1382 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
Xoutput239 net239 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__10583__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ net1449 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_120_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ clknet_leaf_24_wb_clk_i _01783_ _00384_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\]
+ sky130_fd_sc_hd__dfrtp_1
X_06910_ net1123 net895 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07890_ net748 _03830_ net810 vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__o21a_1
X_06841_ net1141 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09560_ _05308_ _05501_ _05190_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a21o_1
XANTENNA__12088__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08894__A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08511_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\]
+ net971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\] net937
+ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o221a_1
X_09491_ _05313_ _05320_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11835__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10929__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08442_ net438 net436 _04382_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__or3_4
XFILLER_0_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07303__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ net935 _04313_ _04314_ net1056 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07324_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\] net727
+ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08464__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09008__A1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07255_ _03193_ _03196_ net820 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout311_A net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07449__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12012__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07186_ net737 _03127_ net1151 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1259_A team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10574__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _06757_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_6
Xfanout1409 net1432 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__clkbuf_4
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_8
XANTENNA_fanout778_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10603__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout433 net434 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 net447 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_8
Xfanout455 _06801_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__buf_6
Xfanout466 net467 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_2
X_09827_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout477 net484 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 _06779_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_8
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_4
XANTENNA_fanout945_A _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ _03243_ _04922_ _05699_ _04818_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12079__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10892__A4 _06403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15160__1541 vssd1 vssd1 vccd1 vccd1 _15160__1541/HI net1541 sky130_fd_sc_hd__conb_1
X_08709_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\] net975
+ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__or2_1
XANTENNA__10629__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11826__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08917__S1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _04537_ net360 _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11434__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ net2024 net301 net341 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07213__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ net2406 _06617_ net350 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__mux2_1
XANTENNA__09131__C net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net2568 net1914 net838 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11054__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07258__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ clknet_leaf_127_wb_clk_i _02134_ _00735_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[724\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11582_ net277 net2760 net455 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ net1279 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
X_10533_ net164 net1029 net1020 net1905 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__A0 _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ net1309 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input74_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ net284 _06277_ net679 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11389__B net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12203_ net1589 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ net1376 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_10395_ net305 net304 _06084_ _06221_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07430__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ net1675 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12065_ _06629_ net2786 net364 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ net494 net646 _06581_ net425 net2040 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14492__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08930__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11817__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ net1390 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
XANTENNA__09486__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12085__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14706_ clknet_leaf_120_wb_clk_i _02470_ _01071_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_11918_ _06619_ net2767 net373 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XANTENNA__08694__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12898_ net1353 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
XANTENNA__08219__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11849_ net276 net2200 net383 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__mux2_1
X_14637_ clknet_leaf_106_wb_clk_i _02401_ _01002_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ clknet_leaf_34_wb_clk_i _02332_ _00933_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08446__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11045__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06962__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13519_ net1278 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XANTENNA__06991__D_N team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14499_ clknet_leaf_25_wb_clk_i _02263_ _00864_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07040_ _02978_ _02981_ net814 vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09097__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11348__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08889__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11899__A3 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\] net1066
+ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07972__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07942_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\] net736
+ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__o221a_1
XANTENNA__10423__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09174__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A2 _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07873_ _03813_ _03814_ net810 vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ net542 _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__nand2_1
X_06824_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] vssd1 vssd1 vccd1 vccd1
+ _02767_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06932__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ net579 _05484_ _05481_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_116_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11284__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ _05085_ _05115_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nor2_1
XANTENNA__11481__C _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11823__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ net1210 _04365_ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout526_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1170_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ net1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\] net967 net919
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07307_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\]
+ net764 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08287_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10795__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14365__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ net1140 _03175_ _03177_ _03178_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__o32a_1
XFILLER_0_14_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout895_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07169_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\]
+ net755 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XANTENNA__12000__A3 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ _06018_ _06019_ _03242_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07963__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11429__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1207 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_8
Xfanout1217 team_03_WB.instance_to_wrap.core.decoder.inst\[16\] vssd1 vssd1 vccd1
+ vccd1 net1217 sky130_fd_sc_hd__buf_4
Xfanout1228 net1229 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1239 team_03_WB.instance_to_wrap.core.decoder.inst\[15\] vssd1 vssd1 vccd1
+ vccd1 net1239 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07208__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 _06546_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_4
Xfanout274 _06446_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
Xfanout285 net286 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07176__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11375__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 _06523_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ clknet_leaf_71_wb_clk_i _01634_ _00235_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09180__A3 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__S1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net1267 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XANTENNA__09468__A1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12752_ net1428 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11391__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11703_ _06745_ net388 net347 net2044 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12683_ net1257 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12784__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14422_ clknet_leaf_93_wb_clk_i _02186_ _00787_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14708__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11634_ _06708_ net389 net354 net2449 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_831 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08428__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14353_ clknet_leaf_97_wb_clk_i _02117_ _00718_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\]
+ sky130_fd_sc_hd__dfrtp_1
X_11565_ net508 net633 _06674_ net488 net2175 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a32o_1
XANTENNA__09640__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ net1291 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
X_10516_ net151 net1029 net1020 net1841 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
X_14284_ clknet_leaf_6_wb_clk_i _02048_ _00649_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\]
+ sky130_fd_sc_hd__dfrtp_1
X_11496_ _06617_ net2739 net396 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__mux2_1
X_13235_ net1264 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10447_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] _06135_ vssd1 vssd1 vccd1
+ vccd1 _06264_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10538__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07817__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ net1283 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
X_10378_ _05986_ _05987_ _06087_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12117_ team_03_WB.instance_to_wrap.WRITE_I _02777_ team_03_WB.instance_to_wrap.wb.curr_state\[0\]
+ _02797_ net2849 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__a32o_1
XANTENNA__11750__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ net1247 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XANTENNA_max_cap324_A _05746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _06617_ net2599 net364 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13999_ clknet_leaf_97_wb_clk_i _01763_ _00364_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11266__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08667__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08210_ net932 _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14388__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07890__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ net441 net433 net589 net553 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__o31a_1
XFILLER_0_111_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11569__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ net1058 net1012 vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09631__A1 _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07300__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07023_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\]
+ net895 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__or3_1
XFILLER_0_114_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10529__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07945__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__B2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[777\]
+ net985 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1016_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold16 team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\] vssd1
+ vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07925_ net1089 net893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\]
+ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__o21a_1
Xhold27 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[2\] vssd1 vssd1 vccd1
+ vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\] vssd1
+ vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 team_03_WB.instance_to_wrap.ADR_I\[29\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout476_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\] net798
+ _03792_ net1113 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06867__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10701__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__A _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07787_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\] net1147
+ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout643_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1385_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net578 _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08658__C1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ _05137_ _05398_ net557 vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout810_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout908_A net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11712__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\]
+ net990 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07881__A0 _03821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _05321_ _05325_ _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__and3_1
XANTENNA__08293__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13755__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08339_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11013__A _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ net507 net630 _06727_ net405 net2057 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__a32o_1
XANTENNA__07633__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] _06142_ vssd1 vssd1
+ vccd1 vccd1 _06143_ sky130_fd_sc_hd__and2_1
X_11281_ net712 _06518_ net824 vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__and3_1
X_13020_ net1350 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10232_ _06071_ _06072_ _03864_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07936__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11193__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ _04862_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] net673 vssd1
+ vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10940__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 net1031 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1036 _05904_ vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_4
XANTENNA_input37_A gpio_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1049 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_14971_ clknet_leaf_40_wb_clk_i _02723_ _01336_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dfrtp_1
X_10094_ _05833_ _05834_ _05841_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__and4_1
Xfanout1058 _02790_ vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__buf_4
XANTENNA__12779__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1069 net1076 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_4
X_13922_ clknet_leaf_129_wb_clk_i _01686_ _00287_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08897__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07372__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08361__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13853_ clknet_leaf_67_wb_clk_i _01617_ _00218_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11248__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ net1311 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14530__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ net713 net701 net303 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__or3b_1
XFILLER_0_97_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13784_ clknet_leaf_11_wb_clk_i _01548_ _00149_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08113__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ net1377 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07872__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12666_ net1370 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07401__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11617_ _06691_ net390 net355 net2381 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
X_14405_ clknet_leaf_108_wb_clk_i _02169_ _00770_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09074__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09613__A1 _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12597_ net1262 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07624__A0 _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11548_ net2499 net489 _06789_ net518 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a22o_1
X_14336_ clknet_leaf_132_wb_clk_i _02100_ _00701_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08821__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold508 team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\] vssd1
+ vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14267_ clknet_leaf_29_wb_clk_i _02031_ _00632_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold519 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\] vssd1
+ vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ net507 net630 _06603_ net400 net2190 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a32o_1
XANTENNA__07547__S net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ net1348 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14198_ clknet_leaf_84_wb_clk_i _01962_ _00563_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11069__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07927__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A2 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ net1375 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1208 team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\] vssd1
+ vssd1 vccd1 vccd1 net2792 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\] vssd1
+ vssd1 vccd1 vccd1 net2803 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\] net1120
+ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__o221a_1
XANTENNA__11487__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08690_ _04626_ _04631_ net869 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08378__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _03578_ _03579_ _03581_ net1117 net1152 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07560__C1 team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06902__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07572_ net1112 _03507_ _03508_ _03510_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__o32a_1
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09213__D _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ net589 _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ _03391_ _05153_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09173_ net439 net431 _05012_ net546 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__o31a_1
XANTENNA__09065__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08124_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\] net789
+ net1011 _04065_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08055_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[246\] net740
+ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o221a_1
XANTENNA__10672__A _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07006_ net606 _02940_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__or3_1
XANTENNA__09238__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08142__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08040__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1300_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\]
+ net987 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\] net925
+ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout760_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\]
+ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__and2_1
XANTENNA__10611__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11478__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ _02948_ _02949_ net529 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__or3b_2
XFILLER_0_93_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08343__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07839_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\]
+ net759 vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11008__A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _06394_ _06447_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nand2_2
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07529__S0 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _05350_ _05366_ net571 vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10781_ _06381_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12520_ net1292 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XANTENNA__07854__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07859__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12451_ net1297 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11402_ net279 net2788 net401 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15170_ net1551 vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08803__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08751__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ net1384 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
X_14121_ clknet_leaf_59_wb_clk_i _01885_ _00486_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11333_ net281 net716 net699 vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14052_ clknet_leaf_20_wb_clk_i _01816_ _00417_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\]
+ sky130_fd_sc_hd__dfrtp_1
X_11264_ net499 net628 _06699_ net414 net2375 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a32o_1
XANTENNA__07909__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ net1254 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XANTENNA__11705__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10215_ _06028_ _06056_ _06026_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a21o_1
X_11195_ net2802 net419 _06678_ net510 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
XANTENNA__08582__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _03109_ _05985_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14954_ clknet_leaf_41_wb_clk_i _02706_ _01319_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dfrtp_1
X_10077_ _03352_ _04475_ net314 vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__mux2_1
XANTENNA__11469__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09531__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ clknet_leaf_94_wb_clk_i _01669_ _00270_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14885_ clknet_leaf_42_wb_clk_i _02648_ _01250_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13920__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13836_ clknet_leaf_8_wb_clk_i _01600_ _00201_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[190\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09611__A _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13767_ clknet_leaf_65_wb_clk_i _01531_ _00132_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\]
+ sky130_fd_sc_hd__dfrtp_1
X_10979_ net266 net2339 net523 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XANTENNA__09834__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__C_N _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12718_ net1341 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13698_ clknet_leaf_131_wb_clk_i _01462_ _00063_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10995__A3 _06569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__D net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ net1256 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14426__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14319_ clknet_leaf_99_wb_clk_i _02083_ _00684_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold305 team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\] vssd1
+ vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07785__B _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 net117 vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold327 team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\] vssd1
+ vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 net178 vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold349 _02607_ vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08248__S1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09860_ _05706_ _05801_ _05718_ _05697_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__or4bb_1
Xfanout807 net811 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10904__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout818 net820 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_4
X_08811_ net1060 _04751_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a21o_1
X_09791_ _05731_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__nor2_1
XANTENNA__10380__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\] vssd1
+ vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\] vssd1
+ vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08742_ _04682_ _04683_ net852 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__o21a_1
Xhold1027 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\] vssd1
+ vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\] vssd1
+ vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\] vssd1
+ vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08325__A1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\] net943
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a221o_1
X_07624_ _03563_ _03565_ net608 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10683__A2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08089__A0 _04029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07555_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\]
+ net777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\] net734
+ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout341_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__A1 _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09825__B2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07836__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ _03425_ _03427_ net608 vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__mux2_2
XFILLER_0_14_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09225_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1289_A team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12882__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1250_A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09589__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1348_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ _05096_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08487__S1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11396__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\]
+ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09087_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\] net933
+ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__o221a_1
XANTENNA__10606__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08800__A2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\]
+ net887 net1037 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__o31a_1
XFILLER_0_130_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold850 team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\] vssd1
+ vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout975_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\] vssd1
+ vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\] vssd1
+ vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold883 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\] vssd1
+ vssd1 vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\] vssd1
+ vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ _05885_ net1810 net287 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09989_ _05874_ net2144 net288 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07772__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10929__D_N team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ net624 _06728_ net463 net369 net1962 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10902_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\] net313 net311 net321
+ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__and4_1
X_14670_ clknet_leaf_58_wb_clk_i _02434_ _01035_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11882_ net643 _06691_ net483 net379 net2078 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13621_ net1430 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ net686 _05517_ _06401_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13552_ net1329 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
X_10764_ net527 _06375_ _06376_ net532 net1717 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14449__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ net1413 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
X_13483_ net1394 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XANTENNA__09029__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10695_ _05583_ _06311_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12434_ net1389 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07055__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15153_ net1534 vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
X_12365_ net1268 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11316_ _06623_ net2818 net411 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__mux2_1
X_14104_ clknet_leaf_12_wb_clk_i _01868_ _00469_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\]
+ sky130_fd_sc_hd__dfrtp_1
X_15084_ net1465 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
X_12296_ net1284 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ clknet_leaf_110_wb_clk_i _01799_ _00400_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ net276 net714 net825 vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10898__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net712 _06517_ _06562_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__or3_1
X_10129_ _05970_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11311__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ clknet_leaf_125_wb_clk_i _02692_ _01302_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11293__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868_ clknet_leaf_54_wb_clk_i net1634 _01233_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08883__C _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__A _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13819_ clknet_leaf_26_wb_clk_i _01583_ _00184_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14799_ clknet_leaf_32_wb_clk_i _02563_ _01164_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07340_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__A2 _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07271_ net1126 _03209_ _03210_ _03212_ net1112 vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a311o_1
X_09010_ net845 _04944_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13816__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15129__1510 vssd1 vssd1 vccd1 vccd1 _15129__1510/HI net1510 sky130_fd_sc_hd__conb_1
XFILLER_0_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11378__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08469__S1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\] vssd1
+ vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold113 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\] vssd1
+ vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net179 vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08794__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\] vssd1
+ vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold146 net211 vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold157 net182 vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13966__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08123__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\] vssd1
+ vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _05706_ _05730_ net324 _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\] vssd1
+ vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout604 _06294_ vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 net618 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08546__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout626 net645 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08546__B2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
X_09843_ _05260_ _05262_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__xnor2_1
Xfanout648 net650 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_4
Xfanout659 _05950_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_2
XANTENNA__08641__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07754__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11484__C _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ _02822_ _02806_ _02801_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__and3b_1
X_09774_ net665 _05715_ _03208_ _04646_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09950__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ net920 _04666_ net1061 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__o21a_1
XANTENNA__07506__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _04596_ _04597_ net853 vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07607_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\]
+ net782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\] net749
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08587_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout723_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _03476_ _03479_ net814 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08077__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11005__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ net1108 _03409_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11720__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ net607 _05147_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nor2_1
X_10480_ net121 net1026 net902 net2469 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07037__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ net584 _05079_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08785__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ net1660 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07993__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _06505_ net2645 net423 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__mux2_1
X_12081_ _06785_ net480 net446 net2127 vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__a22o_1
Xhold680 team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\] vssd1
+ vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10860__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\] vssd1
+ vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ net701 net709 net298 vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__or3b_1
XANTENNA__11541__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ net1415 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14722_ clknet_leaf_118_wb_clk_i _02486_ _01087_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08476__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11934_ net265 net2651 net375 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14653_ clknet_leaf_63_wb_clk_i _02417_ _01018_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_19_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11865_ net297 net2493 net383 vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13604_ net1283 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10816_ _06419_ _06420_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_131_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11796_ net2400 _06626_ net332 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__mux2_1
X_14584_ clknet_leaf_129_wb_clk_i _02348_ _00949_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07276__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13535_ net1273 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
X_10747_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] _05718_ net602 vssd1
+ vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13466_ net1393 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
X_10678_ _02766_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13989__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15205_ net1575 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12021__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net1288 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13397_ net1423 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XANTENNA__07579__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA__09973__A0 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08776__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput218 net218 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_15136_ net1517 vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput229 net229 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12348_ net1355 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XANTENNA__10583__B2 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12279_ net1414 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
X_15067_ net1448 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08528__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ clknet_leaf_130_wb_clk_i _01782_ _00383_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11077__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] vssd1 vssd1 vccd1 vccd1
+ _02783_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10886__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12697__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08510_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\] net920
+ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__o221a_1
XANTENNA__11805__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ _05332_ _05430_ _05315_ _05324_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__o211a_1
XANTENNA__08386__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07503__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14764__CLK clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\] net919
+ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07323_ _03262_ _03264_ net806 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07254_ net803 _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A2 _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08216__B1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\] vssd1
+ vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout304_A _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A0 _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1046_A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__A1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11771__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08519__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _06752_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_6
Xfanout412 _06717_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout423 net424 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_8
Xfanout434 net435 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout467 net485 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
X_09826_ _05764_ _05767_ _05758_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__and3b_2
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout478 net484 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_4
Xfanout489 _06779_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_4
XANTENNA__12079__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _03243_ _04922_ net542 vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout840_A net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06969_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\]
+ net771 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout938_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ net557 _04649_ _04594_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08296__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ net325 _05462_ _05467_ net326 _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08639_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11650_ net2077 _06616_ net350 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ net1699 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] net838 vssd1 vssd1 vccd1
+ vccd1 _02527_ sky130_fd_sc_hd__mux2_1
XANTENNA__07258__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ net278 net2851 net452 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__mux2_1
XANTENNA__11054__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10855__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10532_ net1761 net1029 net1020 team_03_WB.instance_to_wrap.CPU_DAT_I\[7\] vssd1
+ vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ net1279 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10463_ _06134_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ net1263 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XANTENNA__11389__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08044__B _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ net1723 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ net1385 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XANTENNA_input67_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _06080_ _06081_ _06083_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11762__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__C1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12133_ net1700 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07430__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07981__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _06519_ net2748 net363 vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08060__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11514__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14637__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__C1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ net703 _06468_ net822 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10868__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout990 net992 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08930__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13661__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ net1412 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08143__C1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ clknet_leaf_117_wb_clk_i _02469_ _01070_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _06618_ net2652 net376 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08694__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ net1287 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14636_ clknet_leaf_5_wb_clk_i _02400_ _01001_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _06426_ net2045 net381 vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11045__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ clknet_leaf_63_wb_clk_i _02331_ _00932_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\]
+ sky130_fd_sc_hd__dfrtp_1
X_11779_ net2590 _06612_ net332 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10253__A0 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13518_ net1278 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ clknet_leaf_129_wb_clk_i _02262_ _00863_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08235__A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13449_ net1395 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__C net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14167__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__S1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_75_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09410__A2 _04149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15119_ net1500 vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_2
XFILLER_0_76_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08990_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a221o_1
XANTENNA__09066__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07941_ net818 _03876_ net718 vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07872_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\] net748
+ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07185__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ _03280_ _04532_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__or2_1
X_06823_ team_03_WB.instance_to_wrap.core.pc.current_pc\[31\] vssd1 vssd1 vccd1 vccd1
+ _02766_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13316__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__B _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ _05482_ _05483_ net567 vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09005__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ _05413_ _05414_ net556 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
XANTENNA__11284__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11481__D net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10492__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ net1057 _04363_ _04364_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout421_A net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1163_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07306_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\] net727
+ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout519_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08286_ _04224_ _04225_ _04226_ _04227_ net856 net916 vssd1 vssd1 vccd1 vccd1 _04228_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10795__A1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07237_ net1125 _03172_ _03173_ net1131 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1330_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1428_A net1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07984__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07099__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07168_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\]
+ net755 vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout790_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout888_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10614__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[801\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\]
+ net773 net1123 vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07195__S net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07963__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 team_03_WB.instance_to_wrap.core.decoder.inst\[17\] vssd1 vssd1 vccd1
+ vccd1 net1207 sky130_fd_sc_hd__clkbuf_8
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout1229 net1239 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout264 _06537_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
XANTENNA__13684__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _06434_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_2
XANTENNA__08373__C1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 _05946_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09809_ _02923_ _04565_ net665 _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a22o_1
Xfanout297 _06513_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12820_ net1322 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12751_ net1410 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11391__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11702_ _06744_ net389 net346 net2075 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a22o_1
X_12682_ net1257 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ clknet_leaf_87_wb_clk_i _02185_ _00786_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08428__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11633_ _06707_ net391 net354 net2275 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14352_ clknet_leaf_82_wb_clk_i _02116_ _00717_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07597__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11564_ net2067 net488 _06796_ net513 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__a22o_1
XANTENNA__11983__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ net1326 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10515_ net152 net1029 net1020 net1951 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a22o_1
XANTENNA__07651__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11495_ _06616_ net2711 net395 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
X_14283_ clknet_leaf_46_wb_clk_i _02047_ _00648_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09928__A0 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07894__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09585__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13234_ net1422 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
X_10446_ _06032_ _06055_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07939__C1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07403__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _05986_ _05987_ _06087_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__or3_1
X_13165_ net1318 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
X_12116_ _02776_ team_03_WB.instance_to_wrap.READ_I team_03_WB.instance_to_wrap.wb.curr_state\[0\]
+ _02797_ net2868 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a32o_1
X_13096_ net1342 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
X_12047_ _06616_ net2698 net363 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07833__S net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10710__B2 net2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13136__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_122_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12040__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13998_ clknet_leaf_70_wb_clk_i _01762_ _00363_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ net1269 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__08667__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14619_ clknet_leaf_32_wb_clk_i _02383_ _00984_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11018__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07890__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11090__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08140_ net1200 _02820_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09631__A2 _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07642__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ net1183 net876 team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\]
+ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ net1200 _04911_ _04914_ net848 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__o31a_1
XANTENNA__08131__C _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold17 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[6\] vssd1 vssd1 vccd1
+ vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07924_ net613 _03864_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__o21a_2
Xhold28 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[21\] vssd1 vssd1 vccd1
+ vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\] vssd1
+ vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07855_ net1113 _03795_ _03796_ net1127 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13046__A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07786_ _03680_ _03681_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07044__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09525_ _05464_ _05465_ net565 vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08658__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1280_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout636_A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1378_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09456_ net553 _04080_ _04770_ _05135_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06883__A team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08407_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\]
+ net990 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09387_ _05327_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout803_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10609__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08338_ _04274_ _04279_ net868 vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11965__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07094__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11013__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__mux2_1
XANTENNA__07633__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08830__B1 _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] team_03_WB.instance_to_wrap.core.pc.current_pc\[14\]
+ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net516 net640 _06707_ net415 net2117 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10231_ _03864_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11193__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1010 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_2
XFILLER_0_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10940__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1015 _02809_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
Xfanout1026 net1031 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_2
X_14970_ clknet_leaf_31_wb_clk_i _02722_ _01335_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__dfrtp_1
Xfanout1037 _02871_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_8
XFILLER_0_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10093_ net318 _05676_ _05811_ _05931_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__and4bb_1
Xfanout1048 net1049 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08346__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1064 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_4
X_13921_ clknet_leaf_2_wb_clk_i _01685_ _00286_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08897__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08992__S0 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ clknet_leaf_118_wb_clk_i _01616_ _00217_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12803_ net1301 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
X_13783_ clknet_leaf_73_wb_clk_i _01547_ _00148_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ net496 net648 _06569_ net425 net2262 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12734_ net1386 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
XANTENNA__08484__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09614__A1_N team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07872__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15088__1469 vssd1 vssd1 vccd1 vccd1 _15088__1469/HI net1469 sky130_fd_sc_hd__conb_1
X_12665_ net1353 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14404_ clknet_leaf_20_wb_clk_i _02168_ _00769_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\]
+ sky130_fd_sc_hd__dfrtp_1
X_11616_ _06690_ net386 net353 net2369 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09613__A2 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ net1320 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11956__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14335_ clknet_leaf_116_wb_clk_i _02099_ _00700_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\]
+ sky130_fd_sc_hd__dfrtp_1
X_11547_ net641 _06657_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09609__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\] vssd1
+ vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14266_ clknet_leaf_21_wb_clk_i _02030_ _00631_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11971__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08513__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ net2570 net399 _06774_ net513 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10762__B _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13217_ net1265 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
X_10429_ _06248_ _06249_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] net680
+ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14197_ clknet_leaf_89_wb_clk_i _01961_ _00562_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07927__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07129__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13148_ net1351 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13079_ net1417 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
Xhold1209 team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\] vssd1
+ vssd1 vccd1 vccd1 net2793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11487__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11085__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07155__A3 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07640_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\]
+ net760 net1117 vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux4_1
XANTENNA__07560__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ net745 _03511_ _03512_ net1158 vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ net584 _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07312__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10998__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ _05176_ _05182_ _05177_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09172_ _05110_ _05113_ net558 vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09065__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08123_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\]
+ net892 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__or3_1
XANTENNA__11947__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08812__B1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08054_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[86\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\] net727
+ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07005_ _02945_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__and2b_2
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1126_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07039__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08040__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ net941 _04896_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07907_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\]
+ net880 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__and3_1
XANTENNA__11478__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ net568 _04827_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__nor2_2
XANTENNA__07146__A3 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[938\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\]
+ net759 net1117 vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07551__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\] net789
+ _03703_ net1108 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13504__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ net578 _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__or2_1
XANTENNA__07529__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10780_ _06389_ _06380_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and2b_2
XFILLER_0_52_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07502__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07854__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ _05379_ _05380_ net557 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11024__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13872__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07221__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net1364 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11938__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _06413_ net2545 net402 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08803__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ net1382 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09071__A3 _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ clknet_leaf_35_wb_clk_i _01884_ _00485_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07648__S net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ net1038 _06449_ net650 net694 vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__or4_4
XANTENNA__09429__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07082__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14051_ clknet_leaf_19_wb_clk_i _01815_ _00416_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11263_ net1241 net831 _06477_ net668 vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__and4_2
XFILLER_0_123_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11166__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08567__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ net1249 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10214_ _06032_ _06055_ _06030_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__o21ai_1
X_11194_ net654 net706 net267 net697 vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and4_1
X_10145_ _03109_ _05985_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08319__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14953_ clknet_leaf_61_wb_clk_i _02705_ _01318_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dfrtp_1
X_10076_ _05342_ net316 _05919_ net582 _02937_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11469__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13904_ clknet_leaf_83_wb_clk_i _01668_ _00269_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\]
+ sky130_fd_sc_hd__dfrtp_1
X_14884_ clknet_leaf_52_wb_clk_i _02647_ _01249_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10103__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13835_ clknet_leaf_46_wb_clk_i _01599_ _00200_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09611__B _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ clknet_leaf_75_wb_clk_i _01530_ _00131_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09295__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _06551_ _06554_ _06556_ _06391_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__o211a_4
XFILLER_0_58_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07412__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ net1301 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XANTENNA__11641__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ clknet_leaf_2_wb_clk_i _01461_ _00062_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15003__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09047__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12648_ net1351 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
XANTENNA__11929__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_109_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12579_ net1297 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14318_ clknet_leaf_72_wb_clk_i _02082_ _00683_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11944__A3 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\] vssd1
+ vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold317 team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\] vssd1
+ vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold328 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\] vssd1
+ vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold339 team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\] vssd1
+ vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ clknet_leaf_67_wb_clk_i _02013_ _00614_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 net811 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout819 net820 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__buf_4
XANTENNA__11808__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ net1216 _04749_ _04750_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and3_1
XANTENNA__09770__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09770__B2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ _05246_ _05250_ _05269_ net592 vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a31o_1
Xhold1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\] vssd1
+ vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1017 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\] vssd1
+ vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\]
+ net976 team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\] net939
+ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o221a_1
Xhold1028 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\] vssd1
+ vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1039 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\] vssd1
+ vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1390 net1391 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08672_ net924 _04612_ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07533__B1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07623_ _03278_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07554_ _03493_ _03495_ net810 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09825__A2 _05568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07485_ _03426_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__inv_2
XANTENNA__07836__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout334_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09948__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09224_ _05164_ _05165_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ net437 net429 _04267_ net550 vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11396__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1243_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08106_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\]
+ net891 vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__or3_1
XANTENNA__09249__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09086_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\] net918
+ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08037_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\] net788
+ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold840 team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\] vssd1
+ vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold851 team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\] vssd1
+ vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08549__C1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__C _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\] vssd1
+ vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold873 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\] vssd1
+ vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\] vssd1
+ vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11699__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\] vssd1
+ vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_A _04086_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10622__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _05873_ net1844 net288 vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__mux2_1
X_15087__1468 vssd1 vssd1 vccd1 vccd1 _15087__1468/HI net1468 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_95_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10108__C1 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\]
+ net972 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__mux2_1
XANTENNA__08316__A2 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11019__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ net630 _06727_ net468 net372 net2380 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09712__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net316 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[13\]
+ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__o31a_1
X_11881_ net623 _06690_ net463 net377 net2300 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13620_ net1429 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ net275 net2795 net523 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07232__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ net1421 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07288__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ _05798_ net603 vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11623__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net1343 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09029__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10831__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input97_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ net1397 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XANTENNA__08762__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10694_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06316_ net600 vssd1
+ vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14050__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15221_ net912 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12433_ net1304 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15152_ net1533 vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
X_12364_ net1298 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
XANTENNA__08252__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14103_ clknet_leaf_74_wb_clk_i _01867_ _00468_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\]
+ sky130_fd_sc_hd__dfrtp_1
X_11315_ _06622_ net2621 net412 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XANTENNA__07460__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15083_ net1464 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
X_12295_ net1389 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11139__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14034_ clknet_leaf_103_wb_clk_i _01798_ _00399_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\]
+ sky130_fd_sc_hd__dfrtp_1
X_11246_ net503 net621 _06690_ net413 net2294 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a32o_1
XANTENNA__07212__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11177_ net2515 net420 _06668_ net516 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10128_ _05966_ _05967_ _03279_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09504__A1 _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12103__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14936_ clknet_leaf_123_wb_clk_i _02691_ _01301_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10059_ net28 net1033 net907 net2837 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08937__S net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07515__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14867_ clknet_leaf_54_wb_clk_i net1737 _01232_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10768__A _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13818_ clknet_leaf_20_wb_clk_i _01582_ _00183_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\]
+ sky130_fd_sc_hd__dfrtp_1
X_14798_ clknet_leaf_54_wb_clk_i _02562_ _01163_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07142__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07279__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ clknet_leaf_88_wb_clk_i _01513_ _00114_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10822__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\]
+ net898 _03211_ net1149 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__o311a_1
XFILLER_0_128_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08491__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11378__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08779__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08243__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 team_03_WB.instance_to_wrap.core.ru.state\[1\] vssd1 vssd1 vccd1 vccd1 net1687
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold114 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\] vssd1
+ vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold125 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\] vssd1
+ vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\] vssd1
+ vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold147 team_03_WB.instance_to_wrap.ADR_I\[20\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\] vssd1
+ vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _05757_ _05769_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__nand2_1
Xhold169 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[0\] vssd1 vssd1 vccd1
+ vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10950__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08701__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout605 net607 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10889__A0 _06483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout616 net618 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09743__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _05077_ _05783_ _05781_ _05776_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o211a_4
Xfanout627 net629 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_4
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06859__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__A net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ net542 _05713_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__nand2_1
XANTENNA__11484__D net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06985_ net1016 _02814_ _02827_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__or4b_4
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout284_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07601__S0 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08655_ net1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\]
+ net980 team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\] net940
+ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout451_A _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1193_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07606_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08586_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07809__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ net809 _03477_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12893__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1360_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout716_A _06460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07468_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\] net726
+ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o221a_1
XANTENNA__11005__C _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09207_ _03866_ _03947_ _04072_ _05147_ net606 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__a41o_1
XANTENNA__10617__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07399_ net1140 _03338_ _03340_ net1111 vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09138_ _02891_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_1
XANTENNA__12030__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07442__C1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09069_ team_03_WB.instance_to_wrap.core.decoder.inst\[18\] _05010_ _05005_ vssd1
+ vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07993__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ _06626_ net2288 net421 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__mux2_1
X_12080_ _06784_ net483 net446 net2126 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a22o_1
Xhold670 team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\] vssd1
+ vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\] vssd1
+ vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\] vssd1
+ vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ net2207 net428 _06590_ net502 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XANTENNA__11541__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12982_ net1344 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XANTENNA__12097__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ clknet_leaf_125_wb_clk_i _02485_ _01086_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11933_ _06629_ net2662 net375 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ clknet_leaf_127_wb_clk_i _02416_ _01017_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_38_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11864_ net270 net2322 net381 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__mux2_1
XANTENNA__08058__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13603_ net1297 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
X_10815_ net689 _05454_ _06401_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14583_ clknet_leaf_75_wb_clk_i _02347_ _00948_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11795_ net2771 _06625_ net336 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10804__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ net1281 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
X_10746_ net526 _06364_ _06365_ net532 net1689 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08473__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ net1401 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07681__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10677_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06318_ vssd1 vssd1
+ vccd1 vccd1 _06319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08505__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15204_ net912 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ net1378 vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13396_ net1424 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
X_15135_ net1516 vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
X_12347_ net1360 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
Xoutput219 net219 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10583__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15066_ net1447 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12278_ net1343 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
X_14017_ clknet_leaf_0_wb_clk_i _01781_ _00382_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13139__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _06536_ net2488 net492 vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12978__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12088__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09352__A _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11296__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14919_ clknet_leaf_125_wb_clk_i _02674_ _01284_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11835__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08440_ net846 _04368_ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux2_1
XANTENNA__07303__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09498__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07322_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\] net767
+ net736 _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08464__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10945__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15086__1467 vssd1 vssd1 vccd1 vccd1 _15086__1467/HI net1467 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07253_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\] net744
+ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11122__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07184_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\] net754
+ net724 _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08216__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12012__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08134__C _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07424__C1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10574__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__A1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10680__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout402 _06752_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13049__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 net414 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 _06610_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07727__B1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1206_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11523__B2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08924__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net447 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_8
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net460 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_4
X_09825_ _04834_ _05568_ _05765_ net592 _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 net474 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net484 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_2
X_09756_ _05236_ _05661_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__xor2_1
X_06968_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\]
+ net771 vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__mux2_1
XANTENNA__06950__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _04621_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11826__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ _04829_ _05513_ _05627_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout833_A net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06899_ _02837_ net688 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08638_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\] net1204
+ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a221o_1
XANTENNA__10201__A _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11039__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08569_ net851 _04509_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10600_ net2148 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\] net838 vssd1 vssd1 vccd1
+ vccd1 _02528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11580_ net303 net2594 net455 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XANTENNA__10855__B _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07510__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10531_ net2105 net1030 net1020 net2032 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08550__S1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ net1348 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10462_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12201_ net1759 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11211__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ net1366 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] _06142_ vssd1 vssd1
+ vccd1 vccd1 _06220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10871__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07966__B1 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net1602 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10590__B _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ _06628_ net2642 net364 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ net495 net647 _06580_ net425 net2431 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout980 net993 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_4
Xfanout991 net992 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ net1274 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
XANTENNA__11817__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _06617_ net2639 net375 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ clknet_leaf_120_wb_clk_i _02468_ _01069_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10111__A _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12896_ net1378 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ clknet_leaf_38_wb_clk_i _02399_ _01000_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[989\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11847_ _06422_ net2174 net383 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ clknet_leaf_79_wb_clk_i _02330_ _00931_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08446__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11778_ net2623 _06611_ net332 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13517_ net1278 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ net1802 net530 net525 _06356_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14497_ clknet_leaf_0_wb_clk_i _02261_ _00862_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13448_ net1395 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__D _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07406__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ net1424 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ net1499 vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09347__A _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07940_ _03880_ _03881_ net818 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21a_1
X_15049_ net1581 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_44_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08906__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07871_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\] net734
+ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07185__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06822_ net1135 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06932__B2 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _05398_ _05401_ net557 vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09472_ net544 _04296_ _05087_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\]
+ net965 net1067 vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14881__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ net438 net436 _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\]
+ net764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\] net741
+ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07330__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08285_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout414_A _06684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1156_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07236_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\] net794
+ _03171_ net1148 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07167_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1323_A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07098_ net1156 _03038_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout783_A net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1208 net1211 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
Xfanout1219 net1223 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09165__A2 _05106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout950_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout265 _06528_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11726__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net277 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
Xfanout287 net291 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_4
X_09808_ _02923_ _04565_ net543 vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10630__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _06499_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ _03790_ _04953_ _05680_ net665 vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08125__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11027__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ net1341 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07479__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11701_ _06743_ net391 net346 net1998 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12681_ net1252 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XANTENNA__11680__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14420_ clknet_leaf_93_wb_clk_i _02184_ _00785_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08428__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11632_ _06706_ net385 net353 net2745 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ clknet_leaf_98_wb_clk_i _02115_ _00716_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11432__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10077__S net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ net638 net706 _06527_ net697 vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07100__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13302_ net1330 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ net153 net1029 net1020 net1777 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14282_ clknet_leaf_3_wb_clk_i _02046_ _00647_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\]
+ sky130_fd_sc_hd__dfrtp_1
X_11494_ _06615_ net2338 net393 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__mux2_1
XANTENNA__14604__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ net1315 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
X_10445_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] net679 _06260_ _06262_
+ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10538__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__A1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ net1299 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XANTENNA__08061__C1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] _06144_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\]
+ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08071__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ _06287_ _06289_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nand2_1
X_13095_ net1399 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14754__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12046_ _06615_ net2680 net361 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15085__1466 vssd1 vssd1 vccd1 vccd1 _15085__1466/HI net1466 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__B1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ clknet_leaf_110_wb_clk_i _01761_ _00362_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12040__B net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12948_ net1323 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08667__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__S net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ net1407 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
XANTENNA__10776__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13152__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14618_ clknet_leaf_6_wb_clk_i _02382_ _00983_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11423__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14549_ clknet_leaf_92_wb_clk_i _02313_ _00914_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08680__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ net1084 net890 team_03_WB.instance_to_wrap.core.register_file.registers_state\[534\]
+ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14284__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07021_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\] net792
+ net731 _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08278__S0 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11726__A1 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ net941 _04913_ _04912_ net1062 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__o211a_1
X_07923_ _02843_ _03844_ _03863_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\] vssd1
+ vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\] vssd1
+ vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07854_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\] net1158
+ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09016__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__or2_2
XFILLER_0_127_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout364_A _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__inv_2
XANTENNA__08658__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09455_ _05393_ _05396_ net567 vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout531_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06883__B team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout629_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__mux2_1
XANTENNA__13062__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09386_ _04267_ _05326_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08337_ _04275_ _04276_ _04278_ _04277_ net918 net857 vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11965__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08268_ net552 _04179_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11013__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout998_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__o221a_1
XANTENNA__10625__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08199_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__mux2_1
XANTENNA__13651__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10230_ _05012_ net670 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11193__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _06000_ _06001_ _03679_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10940__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1005 net1008 vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1018 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
Xfanout1027 net1031 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__clkbuf_4
X_10092_ _05563_ _05647_ _05933_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand4_1
XANTENNA__07149__A1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08346__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13237__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ clknet_leaf_130_wb_clk_i _01684_ _00285_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08897__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ clknet_leaf_29_wb_clk_i _01615_ _00216_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08992__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14157__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ net1353 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13782_ clknet_leaf_83_wb_clk_i _01546_ _00147_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ net1038 net831 net279 net668 vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__and4_2
XFILLER_0_74_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ net1382 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
XANTENNA__07857__C1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12664_ net1363 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
XANTENNA__08066__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14403_ clknet_leaf_24_wb_clk_i _02167_ _00768_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11615_ _06689_ net390 net354 net2456 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XANTENNA__09074__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09074__B2 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12595_ net1260 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11956__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ clknet_leaf_49_wb_clk_i _02098_ _00699_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07085__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11546_ net520 net634 _06656_ net489 net1766 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10085__A_N _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14265_ clknet_leaf_103_wb_clk_i _02029_ _00630_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\]
+ sky130_fd_sc_hd__dfrtp_1
X_11477_ net638 net706 _06527_ _06558_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12316__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11220__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13216_ net1410 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ net285 _06139_ _06246_ net678 vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__o31a_1
XFILLER_0_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08034__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14196_ clknet_leaf_95_wb_clk_i _01960_ _00561_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ net1360 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
X_10359_ _06191_ _06192_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] net676
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07844__S net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ net1339 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
X_12029_ net624 _06595_ net459 net366 net2355 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07145__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12986__A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07312__A1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10998__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ _04323_ _05179_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09171_ _05111_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09065__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11947__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\] net800
+ net1037 _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__o211a_1
XANTENNA__13610__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08812__A1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08053_ _03992_ _03994_ net807 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07004_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] _02929_ _02827_ _02836_
+ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__or4b_1
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07918__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1021_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A2 _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08955_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\] net986 net925
+ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout481_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\] net778
+ net750 _03847_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08423__S0 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ _04827_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__and2_1
XANTENNA__11883__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1390_A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout746_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08585__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\]
+ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09507_ _05353_ _05374_ net565 vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__mux2_1
XANTENNA__09270__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11635__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _03638_ _03640_ net608 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout913_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09438_ _04593_ _04621_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11024__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ _05310_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ net280 net2838 net401 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XANTENNA__08803__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ net1350 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
X_15084__1465 vssd1 vssd1 vccd1 vccd1 _15084__1465/HI net1465 sky130_fd_sc_hd__conb_1
XFILLER_0_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11331_ _06633_ net2749 net412 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11040__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14050_ clknet_leaf_129_wb_clk_i _01814_ _00415_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\]
+ sky130_fd_sc_hd__dfrtp_1
X_11262_ net494 net615 _06698_ net413 net1982 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11166__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08567__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ net1251 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
X_10213_ _06037_ _06053_ _06035_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11193_ net508 net655 _06677_ net419 net1746 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a32o_1
XANTENNA__08662__S0 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A gpio_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _03109_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08319__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14952_ clknet_leaf_63_wb_clk_i _02704_ _01317_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dfrtp_1
X_10075_ _05346_ _05347_ _05386_ _05341_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09531__A2 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ clknet_leaf_101_wb_clk_i _01667_ _00268_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ clknet_leaf_50_wb_clk_i _02646_ _01248_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11914__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13834_ clknet_leaf_9_wb_clk_i _01598_ _00199_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10429__B2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11626__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13765_ clknet_leaf_108_wb_clk_i _01529_ _00130_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ net691 _06552_ _06553_ _06555_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__a31o_1
XANTENNA__09295__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13697__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12716_ net1298 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
X_13696_ clknet_leaf_132_wb_clk_i _01460_ _00061_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12647_ net1403 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07839__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12578_ net1348 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10601__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ net657 _06641_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__nor2_1
X_14317_ clknet_leaf_106_wb_clk_i _02081_ _00682_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold307 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\] vssd1
+ vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold318 team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\] vssd1
+ vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 net181 vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ clknet_leaf_35_wb_clk_i _02012_ _00613_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08007__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08558__B1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ clknet_leaf_26_wb_clk_i _01943_ _00544_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14322__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout809 net811 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08740_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\] net1001
+ net923 _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__o211a_1
Xhold1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\] vssd1
+ vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\] vssd1
+ vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_03_WB.instance_to_wrap.core.register_file.registers_state\[795\] vssd1
+ vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10117__B1 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1380 net1387 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11865__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1391 net1406 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08671_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\] net1004 net940
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__o221a_1
X_07622_ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] net1016 vssd1 vssd1 vccd1
+ vccd1 _03564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11880__A3 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11617__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\] net777
+ net732 _03494_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07484_ net1155 net1017 net682 vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09223_ _04503_ _05163_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1069_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_840 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09589__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ net437 net429 _04354_ net544 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__o31a_1
XANTENNA__08246__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08105_ _04045_ _04046_ net813 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11396__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09085_ _05021_ _05026_ net868 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1236_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08036_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\]
+ net887 net1011 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__o31a_1
XFILLER_0_128_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput90 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold830 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\] vssd1
+ vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 net192 vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\] vssd1
+ vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold863 team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\] vssd1
+ vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold874 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\] vssd1
+ vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold885 team_03_WB.instance_to_wrap.ADR_I\[26\] vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1403_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold896 team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\] vssd1
+ vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09265__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _05872_ net1786 net287 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout863_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07772__A1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net1213 _04879_ _04878_ net1206 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11856__A0 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11019__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _04770_ _04809_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ net691 _05659_ net587 vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11880_ net641 _06689_ net481 net380 net2291 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a32o_1
XANTENNA__09712__B _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _06431_ _06433_ _06401_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11035__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ net1429 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07288__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ _02775_ _06294_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ net1260 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13481_ net1397 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XANTENNA__09029__A1 net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ net1633 net531 net526 _06332_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15220_ net1580 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_12432_ net1417 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__12033__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08344__A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15151_ net1532 vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
X_12363_ net1253 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10595__B1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14102_ clknet_leaf_86_wb_clk_i _01866_ _00467_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\]
+ sky130_fd_sc_hd__dfrtp_1
X_11314_ _06479_ net2769 net410 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__mux2_1
X_15082_ net1463 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_121_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07460__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ net1411 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XANTENNA__11139__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11909__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14033_ clknet_leaf_94_wb_clk_i _01797_ _00398_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[387\]
+ sky130_fd_sc_hd__dfrtp_1
X_11245_ net1242 net832 net278 net668 vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07394__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ net640 _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07763__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__A0 _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09504__A2 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14935_ clknet_leaf_125_wb_clk_i _02690_ _01300_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10058_ net29 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1
+ vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07515__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08712__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11644__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14866_ clknet_leaf_54_wb_clk_i net2718 _01231_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10768__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07423__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817_ clknet_leaf_112_wb_clk_i _01581_ _00182_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14797_ clknet_leaf_32_wb_clk_i _02561_ _01162_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07279__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08953__S net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13748_ clknet_leaf_91_wb_clk_i _01512_ _00113_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13679_ clknet_leaf_100_wb_clk_i _01443_ _00044_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12024__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11378__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08779__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10586__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\] vssd1
+ vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold115 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[28\] vssd1 vssd1 vccd1
+ vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold126 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[20\] vssd1 vssd1 vccd1
+ vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\] vssd1
+ vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _02623_ vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold159 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\] vssd1
+ vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ net317 _05851_ _05429_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__or3b_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_2
X_09841_ _02992_ _05671_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__o21ai_1
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08400__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 net629 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__buf_2
XANTENNA__07754__A1 net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 net644 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09772_ net540 _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_1
X_06984_ _02828_ _02829_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__or3_2
X_08723_ net937 _04664_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11838__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A _06430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15083__1464 vssd1 vssd1 vccd1 vccd1 _15083__1464/HI net1464 sky130_fd_sc_hd__conb_1
X_08654_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\] net1004
+ net924 _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10510__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07601__S1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\]
+ net881 vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__and3_1
XANTENNA__14218__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout444_A net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1186_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07536_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\] net731
+ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08467__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07467_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\] net739
+ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11005__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1353_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _03866_ _04072_ _05147_ net606 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a31o_1
XANTENNA__12015__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07690__B1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07398_ net1121 _03335_ _03339_ net1131 vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09137_ net529 _02944_ _02948_ _02952_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10577__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09068_ net1062 _05009_ _05008_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__a21o_1
XANTENNA__07442__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout980_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07993__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ net1157 _03953_ _03952_ net1140 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o211a_1
XANTENNA__10633__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold660 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\] vssd1
+ vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold671 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\] vssd1
+ vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10860__C net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold682 team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\] vssd1
+ vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net621 _06589_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__nor2_1
Xhold693 team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\] vssd1
+ vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07745__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08942__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12981_ net1263 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XANTENNA__11829__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10869__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ clknet_leaf_125_wb_clk_i _02484_ _01085_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11932_ _06519_ net2631 net376 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14651_ clknet_leaf_30_wb_clk_i _02415_ _01016_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\]
+ sky130_fd_sc_hd__dfstp_1
X_11863_ _06682_ net469 net382 net2030 vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13602_ net1283 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
X_10814_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[27\] _05865_ net321 _06403_
+ net687 vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a41o_1
X_11794_ net2723 _06624_ net336 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__mux2_1
X_14582_ clknet_leaf_92_wb_clk_i _02346_ _00947_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_71_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10804__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _05706_ net602 vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__nand2_1
X_13533_ net1273 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12006__A0 _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13464_ net1395 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XANTENNA__07681__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] _06317_ vssd1 vssd1
+ vccd1 vccd1 _06318_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15203_ net911 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12415_ net1374 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13395_ net1421 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09422__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07028__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10568__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12021__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07433__B1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12346_ net1372 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
X_15134_ net1515 vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_121_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08630__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_116_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15065_ net1446 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_121_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12277_ net1267 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XANTENNA__13885__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14016_ clknet_leaf_134_wb_clk_i _01780_ _00381_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\]
+ sky130_fd_sc_hd__dfrtp_1
X_11228_ net269 net2408 net492 vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XANTENNA__09725__A2 _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11159_ net1040 net834 net300 net667 vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13155__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11296__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14918_ clknet_leaf_125_wb_clk_i _02673_ _01283_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08249__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__C_N net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14849_ clknet_leaf_54_wb_clk_i net1609 _01214_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11048__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ _04310_ _04311_ net1210 vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__o21a_1
XANTENNA__08449__C1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08683__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06992__A _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07321_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\]
+ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07252_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\] net732
+ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11122__B net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07183_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\] net787
+ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__or2_1
XANTENNA__10559__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08134__D _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10961__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11776__C net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout403 _06752_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_6
Xfanout414 _06684_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_4
Xfanout425 net428 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout436 _04079_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11523__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_A _06778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08924__B1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout447 _06819_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__buf_4
X_09824_ _05073_ _05688_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout458 net460 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1101_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 net471 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__14040__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06967_ net1157 _02907_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__and3_1
X_09755_ net583 _05276_ _05687_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a31o_2
XANTENNA__10689__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06950__A2 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08706_ net441 net433 _04647_ net547 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__o31a_1
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09686_ _03988_ _04178_ _04820_ _03985_ net1018 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__a32o_1
XANTENNA__08159__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06898_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] _02815_ _02828_
+ _02831_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__or4_1
XFILLER_0_59_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08637_ _04573_ _04578_ net869 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout826_A _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14190__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11039__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08568_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\] net934
+ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07519_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[870\] net1148
+ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__a221o_1
X_08499_ net1062 _04438_ _04439_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__or3_1
XANTENNA__10628__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09652__B2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10530_ net167 net1030 net1021 net1884 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08860__C1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11032__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ _06043_ _06050_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12200_ net1716 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13180_ net1352 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10392_ _06218_ _06219_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] net677
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08612__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10871__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07966__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11762__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net1678 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10970__B1 _06549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ _06627_ net2754 net362 vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold490 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\] vssd1
+ vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07718__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _06453_ net703 net822 vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10722__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout970 net993 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_4
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout992 net993 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__buf_2
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ net1306 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
XANTENNA__14533__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\] vssd1
+ vssd1 vccd1 vccd1 net2774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ clknet_leaf_11_wb_clk_i _02467_ _01068_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11915_ _06616_ net2725 net375 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ net1376 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11922__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ clknet_leaf_2_wb_clk_i _02398_ _00999_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\]
+ sky130_fd_sc_hd__dfstp_1
X_11846_ net279 net2277 net381 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ clknet_leaf_123_wb_clk_i _02329_ _00930_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\]
+ sky130_fd_sc_hd__dfrtp_1
X_11777_ net2452 _06609_ net335 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10728_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] _05632_ net601 vssd1
+ vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__mux2_1
X_13516_ net1278 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14496_ clknet_leaf_134_wb_clk_i _02260_ _00861_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ net1396 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
X_10659_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\] team_03_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ net840 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15082__1463 vssd1 vssd1 vccd1 vccd1 _15082__1463/HI net1463 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07406__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ net1421 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XANTENNA__07957__A1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ net1498 vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_2
XFILLER_0_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ net1247 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15048_ net135 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14063__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07709__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _03808_ _03811_ net819 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09174__A3 _05068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ _05394_ _05400_ net564 vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_13_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09471_ net552 _04149_ _05090_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_56_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10021__B net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__C1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08422_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\]
+ net965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\] net1202
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10956__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07304_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\]
+ net892 vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07645__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11441__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07235_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\] net794
+ net747 _03176_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1149_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07166_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] net1012 _03107_ vssd1
+ vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07984__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08442__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14406__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11744__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07097_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[993\] net1123
+ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1316_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09972__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15178__1559 vssd1 vssd1 vccd1 vccd1 _15178__1559/HI net1559 sky130_fd_sc_hd__conb_1
XANTENNA__12899__A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1211 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08373__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _06557_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_2
XANTENNA__09273__A _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _06430_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_2
X_09807_ _05268_ _05747_ _05748_ net592 vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a211oi_2
Xfanout288 net290 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_4
X_07999_ net808 _03939_ _03940_ net815 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__o211a_1
Xfanout299 _06495_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__buf_2
XANTENNA_fanout943_A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09738_ net543 _05679_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08125__A1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11027__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net591 _05598_ _05599_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__o31ai_4
XANTENNA__09873__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11742__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09873__B2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11700_ _06742_ net389 net346 net1833 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__a22o_1
X_12680_ net1292 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11631_ _06705_ net389 net354 net2586 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09086__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11043__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14350_ clknet_leaf_70_wb_clk_i _02114_ _00715_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11432__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ net2073 net488 _06795_ net513 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10513_ net2567 net1023 net1019 net2134 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
X_13301_ net1330 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ clknet_leaf_67_wb_clk_i _02045_ _00646_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11493_ _06614_ net2779 net395 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13232_ net1429 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
XANTENNA_input72_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ net284 _06136_ _06261_ net679 vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__o31ai_1
XANTENNA__09448__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07939__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13163_ net1276 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
X_10375_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] net677 _06203_ _06205_
+ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__A3 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12114_ net1134 net1973 _06292_ net1137 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13094_ net1427 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11917__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ _06614_ net2655 net363 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13996_ clknet_leaf_5_wb_clk_i _01760_ _00361_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12040__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09911__A _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ net1265 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
XANTENNA__07324__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09864__B2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11652__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ net1337 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09122__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ clknet_leaf_104_wb_clk_i _02381_ _00982_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _06663_ net462 net331 net2343 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08824__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ clknet_leaf_92_wb_clk_i _02312_ _00913_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14429__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_131_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14479_ clknet_leaf_99_wb_clk_i _02243_ _00844_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10792__A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07020_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\]
+ net895 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08278__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11187__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08052__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09792__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08971_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07922_ net1229 net1012 _03107_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09001__C1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\] vssd1
+ vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[955\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[923\]
+ net781 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__mux2_1
XANTENNA__07606__A net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07563__C1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _03700_ _03701_ _03722_ net614 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__o211a_2
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ _05372_ _05376_ net563 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11111__A0 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1099_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__D_N _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _05394_ _05395_ net557 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10465__A2 net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09032__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08405_ net1200 _04343_ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09385_ _04267_ _05326_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__nor2_1
XANTENNA__10870__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout524_A _06395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1266_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07618__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08815__C1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ net439 net431 _04207_ net546 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__o31a_1
XANTENNA__07094__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\] net1116
+ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08198_ net929 _04138_ _04139_ net850 vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07149_ net804 _03086_ _03089_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07397__A2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ _03679_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nor3_1
XFILLER_0_112_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13946__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1006 net1008 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11737__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10091_ _05583_ _05596_ _05821_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__and4b_1
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
XANTENNA__10641__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1028 net1031 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08346__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1039 _02793_ vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11350__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11038__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13850_ clknet_leaf_22_wb_clk_i _01614_ _00215_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12801_ net1287 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XANTENNA__09731__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15081__1462 vssd1 vssd1 vccd1 vccd1 _15081__1462/HI net1462 sky130_fd_sc_hd__conb_1
X_10993_ net2656 net425 _06568_ net504 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
X_13781_ clknet_leaf_89_wb_clk_i _01545_ _00146_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[135\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07306__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13253__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12732_ net1346 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12663_ net1413 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
X_14402_ clknet_leaf_131_wb_clk_i _02166_ _00767_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\]
+ sky130_fd_sc_hd__dfrtp_1
X_11614_ _06688_ net385 net353 net2593 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12594_ net1419 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ clknet_leaf_76_wb_clk_i _02097_ _00698_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ net2132 net486 _06788_ net500 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XANTENNA__08821__A2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14264_ clknet_leaf_9_wb_clk_i _02028_ _00629_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\]
+ sky130_fd_sc_hd__dfrtp_1
X_11476_ net2546 net400 _06773_ net517 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11708__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ net305 net304 _06063_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__a211o_1
XANTENNA__11220__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ net1378 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14195_ clknet_leaf_113_wb_clk_i _01959_ _00560_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10916__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ net283 _06148_ _06186_ net676 vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o31a_1
XANTENNA__09906__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ net1366 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08810__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__C1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11647__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13077_ net1268 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
X_10289_ _05963_ _06128_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06869__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07426__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ _06770_ net476 net367 net2598 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13979_ clknet_leaf_30_wb_clk_i _01743_ _00344_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06984__B _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07848__A0 _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11644__A1 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15177__1558 vssd1 vssd1 vccd1 vccd1 _15177__1558/HI net1558 sky130_fd_sc_hd__conb_1
XFILLER_0_111_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09170_ net443 net435 _04922_ net547 vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08691__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09696__S0 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08121_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\]
+ net891 vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07076__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09470__C1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\] net767
+ net728 _03993_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13969__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ _02838_ _02928_ _02935_ _02832_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__o211a_2
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__C1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__A0 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07784__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13338__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07336__A team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\]
+ net881 vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__and3_1
X_08885_ net549 _04825_ _04772_ net564 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__a211o_1
XANTENNA__08423__S1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout474_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07536__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\] net1117
+ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07551__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout641_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\]
+ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1383_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _04778_ _05441_ _05444_ _05446_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_17_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07698_ net682 _03639_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and2b_1
XANTENNA__08500__A1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ _04566_ _04680_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_133_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11024__C net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ _05176_ _05181_ _05309_ _05177_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__o211a_1
XANTENNA__11399__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\] net928
+ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09299_ _04619_ _05238_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__and2_1
XANTENNA__10636__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11330_ _06632_ net2575 net411 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11040__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ net710 net273 net822 vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08567__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10212_ _06037_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nand2_1
X_13000_ net1340 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11192_ net1040 net833 _06545_ net667 vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__and4_1
XANTENNA__10374__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _04148_ net670 _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08319__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14951_ clknet_leaf_40_wb_clk_i _02703_ _01316_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input35_A gpio_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11323__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ clknet_leaf_72_wb_clk_i _01666_ _00267_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\]
+ sky130_fd_sc_hd__dfrtp_1
X_14882_ clknet_leaf_52_wb_clk_i _02645_ _01247_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_13833_ clknet_leaf_48_wb_clk_i _01597_ _00198_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13764_ clknet_leaf_8_wb_clk_i _01528_ _00129_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10976_ net691 _05142_ _02932_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ net1254 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13695_ clknet_leaf_121_wb_clk_i _01459_ _00060_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11930__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12646_ net1423 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08805__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ net1287 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10062__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ clknet_leaf_8_wb_clk_i _02080_ _00681_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\]
+ sky130_fd_sc_hd__dfrtp_1
X_11528_ net497 net620 _06640_ net486 net1848 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\] vssd1
+ vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 net228 vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14247_ clknet_leaf_65_wb_clk_i _02011_ _00612_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ net2498 net398 _06766_ net499 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08102__S0 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14178_ clknet_leaf_126_wb_clk_i _01942_ _00543_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[532\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13129_ net1251 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1008 team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\] vssd1
+ vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11314__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1019 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\] vssd1
+ vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12997__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14617__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1370 net1372 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__buf_4
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08670_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__mux2_1
Xfanout1381 net1383 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__buf_4
XANTENNA__08686__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1392 net1394 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__buf_4
XANTENNA__09371__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ net722 _03562_ _03546_ _03538_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07552_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\]
+ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__and2_1
XANTENNA__14767__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12001__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07297__A1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07483_ _03407_ _03408_ _03416_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o22a_2
XFILLER_0_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09222_ _04503_ _05163_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09153_ net550 _04384_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08104_ net1108 _04042_ _04043_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__or3_1
XANTENNA__11141__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06880__D team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ net1210 _05024_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08035_ _03974_ _03976_ net1157 vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__o21ai_1
Xhold820 team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\] vssd1
+ vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xinput80 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15080__1461 vssd1 vssd1 vccd1 vccd1 _15080__1461/HI net1461 sky130_fd_sc_hd__conb_1
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput91 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_1
XFILLER_0_25_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1131_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08549__A1 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\] vssd1
+ vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold842 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\] vssd1
+ vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold853 team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\] vssd1
+ vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold864 team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\] vssd1
+ vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\] vssd1
+ vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold886 _02629_ vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\] vssd1
+ vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ _05871_ net1903 net290 vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__mux2_1
XANTENNA__09980__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14297__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10108__A1 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\]
+ net972 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout856_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ _02937_ net549 net559 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\] net786
+ net725 _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o211a_1
X_08799_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[33\] net976
+ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10830_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[24\] net307 _06432_ net690
+ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07288__A1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__B _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net527 _06373_ _06374_ net532 net2135 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a32o_1
XANTENNA__07232__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12500_ net1320 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_10692_ net600 _06313_ _06329_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a31oi_2
X_13480_ net1397 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
X_12431_ net1407 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08332__S0 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11051__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ net1531 vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net1248 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07996__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14101_ clknet_leaf_88_wb_clk_i _01865_ _00466_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07460__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _06621_ net2696 net409 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux2_1
X_15081_ net1462 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ net1287 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11244_ net518 net641 _06689_ net415 net2098 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a32o_1
X_14032_ clknet_leaf_83_wb_clk_i _01796_ _00397_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08360__A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07212__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net694 net713 net297 vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__or3b_1
X_15176__1557 vssd1 vssd1 vccd1 vccd1 _15176__1557/HI net1557 sky130_fd_sc_hd__conb_1
X_10126_ _03279_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07763__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08960__A1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06971__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net30 net1032 net906 net2861 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__o22a_1
X_14934_ clknet_leaf_126_wb_clk_i _02689_ _01299_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08173__C1 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ clknet_leaf_53_wb_clk_i net2470 _01230_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10093__B_N _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13816_ clknet_leaf_11_wb_clk_i _01580_ _00181_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14796_ clknet_leaf_62_wb_clk_i _02560_ _01161_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07279__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07142__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ clknet_leaf_112_wb_clk_i _01511_ _00112_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _06538_ _06539_ _06540_ _06399_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o211a_4
XANTENNA__11660__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13678_ clknet_leaf_70_wb_clk_i _01442_ _00043_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08535__A _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08228__B1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ net1262 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XANTENNA__09425__C1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__A0 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10035__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__B2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07987__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 team_03_WB.instance_to_wrap.ADR_I\[9\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold116 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\] vssd1
+ vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold127 _02519_ vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[1\] vssd1 vssd1 vccd1
+ vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\] vssd1
+ vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08270__A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09840_ net574 _05447_ _05439_ net580 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a211o_1
Xfanout607 _02938_ vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08400__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout618 net626 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout629 net645 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__buf_2
XFILLER_0_123_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08951__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ _03208_ _04646_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06983_ _02806_ _02810_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13616__A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12520__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08653_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\] net979
+ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07604_ net819 _03545_ net722 vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__a21o_1
X_08584_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\]
+ net795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\] net746
+ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1081_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__A3 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10813__A2 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ net817 _03401_ net717 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ net529 _03491_ _04074_ _05144_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and4_2
XFILLER_0_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09416__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\] net791
+ _03334_ net1146 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout604_A _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1346_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09975__S net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ net584 _05076_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nand2_1
XANTENNA__10577__B2 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\]
+ net991 net926 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__mux4_1
XANTENNA__07442__A1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08018_ net728 _03957_ _03959_ net1152 vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__a211o_1
Xhold650 team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\] vssd1
+ vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold661 net188 vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout973_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\] vssd1
+ vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\] vssd1
+ vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10860__D _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold694 team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\] vssd1
+ vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13687__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__A3 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _03241_ net661 vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09723__B _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ net1322 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__B _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _06628_ net2595 net376 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11046__A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14650_ clknet_leaf_6_wb_clk_i _02414_ _01015_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\]
+ sky130_fd_sc_hd__dfstp_1
X_11862_ net298 net1975 net384 vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13601_ net1278 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
X_10813_ _05866_ net320 _06404_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__o31a_1
XFILLER_0_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14581_ clknet_leaf_87_wb_clk_i _02345_ _00946_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\]
+ sky130_fd_sc_hd__dfstp_1
X_11793_ net2798 _06623_ net333 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ net1273 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] net602 vssd1 vssd1 vccd1
+ vccd1 _06364_ sky130_fd_sc_hd__or2_1
XANTENNA__10804__A2 _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13463_ net1395 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07681__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10675_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06316_ vssd1 vssd1
+ vccd1 vccd1 _06317_ sky130_fd_sc_hd__or2_1
XANTENNA__09958__A0 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ net911 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12414_ net1384 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XANTENNA__08505__D _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13394_ net1329 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11765__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ net1514 vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
X_12345_ net1356 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08630__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ net1445 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
X_12276_ net1323 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11517__A0 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14015_ clknet_leaf_114_wb_clk_i _01779_ _00380_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\]
+ sky130_fd_sc_hd__dfrtp_1
X_11227_ _06527_ net2330 net492 vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XANTENNA__10125__A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08394__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ net520 net657 _06656_ net420 net1825 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a32o_1
XANTENNA__10740__A1 _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11655__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ _04770_ net672 _05949_ _03060_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11089_ _06621_ net2755 net421 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08146__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07434__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14917_ clknet_leaf_125_wb_clk_i _02672_ _01282_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11296__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ clknet_leaf_54_wb_clk_i net1690 _01213_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11048__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ clknet_leaf_60_wb_clk_i _02543_ _01144_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07320_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\] net764
+ net740 _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a211o_1
XANTENNA__13171__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07251_ _03190_ _03192_ net808 vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07672__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10008__A0 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07182_ net1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\]
+ net754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\] net737
+ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11122__C net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11756__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07424__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11771__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout404 _06752_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_4
Xfanout415 net416 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08924__A1 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout437 net438 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_2
X_09823_ _05265_ _05267_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09824__A _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_8
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ net358 _05569_ _05690_ _05691_ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__a221o_1
X_06966_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\] net1122
+ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a221o_1
XANTENNA__09035__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08705_ _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__inv_2
X_09685_ net663 _05626_ _03988_ _04178_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_55_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout554_A _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06897_ _02815_ _02828_ _02832_ _02794_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and4bb_1
XANTENNA_fanout1296_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08636_ net1060 _04576_ _04577_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07360__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11039__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\] net919
+ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout721_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_54_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13081__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07518_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] net821 vssd1 vssd1 vccd1
+ vccd1 _03460_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08498_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\]
+ net989 net1075 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__mux4_1
XANTENNA__07112__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09652__A2 _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15175__1556 vssd1 vssd1 vccd1 vccd1 _15175__1556/HI net1556 sky130_fd_sc_hd__conb_1
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11995__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ _03389_ _03390_ net608 vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__mux2_4
XFILLER_0_130_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08860__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ net305 net304 _06043_ _06050_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08903__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11747__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07415__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10391_ net283 _06144_ _06215_ net681 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o31a_1
XANTENNA__10644__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ net1669 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _06505_ net2516 net363 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__mux2_1
Xhold480 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\] vssd1
+ vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold491 team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\] vssd1
+ vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012_ net502 net651 _06579_ net428 net2002 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__clkbuf_4
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__clkbuf_4
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 _04086_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07254__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12963_ net1297 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\] vssd1
+ vssd1 vccd1 vccd1 net2764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14702_ clknet_leaf_39_wb_clk_i _02466_ _01067_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.SEL_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\] vssd1
+ vssd1 vccd1 vccd1 net2775 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _06615_ net2681 net373 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12894_ net1381 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14633_ clknet_leaf_60_wb_clk_i _02397_ _00998_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__14828__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11845_ _06413_ net2116 net384 vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14564_ clknet_leaf_16_wb_clk_i _02328_ _00929_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ net1039 _06462_ net387 vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__and3_1
XANTENNA__08300__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__A0 _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ net1278 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10727_ net1850 net533 net528 _06355_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a22o_1
XANTENNA__08851__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14495_ clknet_leaf_109_wb_clk_i _02259_ _00860_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13852__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13446_ net1401 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10658_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ net840 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07406__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ net1329 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10589_ net1134 team_03_WB.instance_to_wrap.WRITE_I net1137 _06292_ vssd1 vssd1 vccd1
+ vccd1 _02534_ sky130_fd_sc_hd__a22o_1
XANTENNA__12335__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15116_ net1497 vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12328_ net1285 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09159__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
X_12259_ net1297 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08906__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06917__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08119__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09470_ net570 _05407_ _05411_ net326 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__o211a_1
XFILLER_0_91_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07342__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08421_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\]
+ net965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\] net1068
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07893__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ _04280_ _04293_ net844 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_4
XFILLER_0_47_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11977__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07645__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11441__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08283_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[727\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07234_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or3_1
XANTENNA__06942__S net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08723__A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07165_ _02808_ net1013 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1
+ vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o21a_4
XFILLER_0_131_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout302_A _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08442__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1044_A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07096_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[865\]
+ net876 _03037_ net1150 vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__a311o_1
XFILLER_0_30_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1309_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09554__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout671_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout267 _06550_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07030__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _05268_ _05747_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 _06426_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_2
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_2
X_07998_ _03935_ _03936_ net808 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07581__B1 _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _03790_ _04953_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__or2_1
X_06949_ net609 _02888_ _02890_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout936_A _04087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ net326 _05533_ _05603_ net359 _05608_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a221oi_4
XANTENNA__11027__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08619_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\]
+ net970 net1071 vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux4_1
XANTENNA__10639__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ net591 _05519_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__o21a_1
XANTENNA__11680__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11630_ _06704_ net386 net353 net2286 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XANTENNA__09086__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07097__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11432__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ net655 _06671_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13300_ net1393 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10640__A0 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ net2180 net1028 net1022 net2072 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14280_ clknet_leaf_27_wb_clk_i _02044_ _00645_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11492_ _06613_ net2824 net393 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ net1388 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
X_10443_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] _06135_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08597__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07249__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08061__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input65_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ net1256 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10374_ net286 _06204_ net677 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08071__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ net1135 net1973 _06282_ team_03_WB.instance_to_wrap.core.ru.state\[5\] vssd1
+ vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13093_ net1274 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
X_12044_ _06613_ net2848 net361 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout790 net796 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13995_ clknet_leaf_17_wb_clk_i _01759_ _00360_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14650__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11933__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ net1398 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07324__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08521__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12877_ net1290 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11234__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14616_ clknet_leaf_10_wb_clk_i _02380_ _00981_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[970\]
+ sky130_fd_sc_hd__dfstp_1
X_11828_ _06661_ net461 net331 net1934 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a22o_1
XANTENNA__09077__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07627__A1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14547_ clknet_leaf_115_wb_clk_i _02311_ _00912_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11759_ net657 _06585_ net472 net339 net2167 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a32o_1
XANTENNA__08824__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10631__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14478_ clknet_leaf_70_wb_clk_i _02242_ _00843_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13429_ net1313 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11187__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_100_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08970_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\]
+ net1008 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\] net925
+ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07921_ net1132 _03852_ _03862_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13748__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07852_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\] net734
+ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__o221a_1
X_15174__1555 vssd1 vssd1 vccd1 vccd1 _15174__1555/HI net1555 sky130_fd_sc_hd__conb_1
XFILLER_0_39_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_2
X_07783_ net610 _03724_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__nor2_1
XANTENNA__11843__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13624__A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _05351_ _05373_ net562 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13898__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06937__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07622__A team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _05109_ _05112_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__nor2_1
XANTENNA__10459__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08404_ net943 _04345_ _04344_ net1062 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__o211a_1
XANTENNA__11144__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09384_ _03529_ _05157_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08335_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08815__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__A2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1161_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ net439 net431 _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__nor3_1
XANTENNA__11965__A3 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08830__A3 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07217_ net1151 _03158_ _03155_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21a_1
X_08197_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\] net913
+ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout1426_A net1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09983__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08043__A1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ net749 _03088_ net809 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_A net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07079_ _03016_ _03020_ _03019_ net1111 vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09284__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1007 net1008 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__clkbuf_2
X_10090_ _05623_ _05632_ _05659_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1018 _02803_ vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__clkbuf_4
Xfanout1029 net1030 vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11350__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ net1379 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ clknet_leaf_91_wb_clk_i _01544_ _00145_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07306__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ net625 _06567_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07532__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ net1361 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XANTENNA__07857__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09059__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12662_ net1346 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14401_ clknet_leaf_0_wb_clk_i _02165_ _00766_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08066__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11613_ _06687_ net386 net353 net2205 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08806__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ net1311 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ clknet_leaf_128_wb_clk_i _02096_ _00697_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[686\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07085__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11956__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net649 _06654_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14263_ clknet_leaf_75_wb_clk_i _02027_ _00628_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07490__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11475_ net656 _06600_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11169__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13214_ net1386 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
X_10426_ _06021_ _06062_ _06017_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08034__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14194_ clknet_leaf_105_wb_clk_i _01958_ _00559_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10916__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09782__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11928__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ net1357 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
X_10357_ net283 _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nand2_1
XANTENNA__09906__B _05833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10832__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12613__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07793__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08990__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07707__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ net1322 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
X_10288_ _05363_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12027_ _06769_ net462 net365 net2549 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07545__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A2 _06701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__S0 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13978_ clknet_leaf_23_wb_clk_i _01742_ _00343_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12929_ net1289 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10852__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08120_ _04059_ _04061_ net1154 vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__o21a_1
XANTENNA__09696__S1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08051_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\]
+ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07002_ net605 _02940_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_128_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08025__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10742__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08953_ _04863_ _04894_ net554 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07904_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\] net732
+ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07336__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ net547 _04825_ _04772_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07536__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__C1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07835_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout467_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07766_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11096__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14076__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _04416_ _04446_ _04505_ _04533_ net551 net562 vssd1 vssd1 vccd1 vccd1 _05447_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07352__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11635__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] net1016 vssd1 vssd1 vccd1
+ vccd1 _03639_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1376_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__S net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09436_ _05374_ _05377_ net566 vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07814__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ _05183_ _05190_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or3_1
XFILLER_0_35_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout801_A _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11024__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07498__S net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ net1071 _04258_ _04259_ net870 vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o31a_1
XANTENNA__09279__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08264__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07472__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net1055 _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ net494 net615 _06697_ net413 net2228 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a32o_1
XFILLER_0_133_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10211_ _06051_ _06052_ _06040_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__a21o_1
XANTENNA__09764__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11191_ net2158 net419 _06676_ net510 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11571__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__C1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] net670 vssd1 vssd1 vccd1
+ vccd1 _05984_ sky130_fd_sc_hd__nand2_1
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11049__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14950_ clknet_leaf_61_wb_clk_i _02702_ _01315_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10073_ _02814_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__or2_1
X_13901_ clknet_leaf_104_wb_clk_i _01665_ _00266_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\]
+ sky130_fd_sc_hd__dfrtp_1
X_14881_ clknet_leaf_50_wb_clk_i _02644_ _01246_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13832_ clknet_leaf_18_wb_clk_i _01596_ _00197_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09819__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11087__A0 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ clknet_leaf_25_wb_clk_i _01527_ _00128_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11626__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10975_ _02829_ net690 _06552_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14569__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12714_ net1249 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ clknet_leaf_48_wb_clk_i _01458_ _00059_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ net1275 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XANTENNA__10827__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08093__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ net1408 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15173__1554 vssd1 vssd1 vccd1 vccd1 _15173__1554/HI net1554 sky130_fd_sc_hd__conb_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14315_ clknet_leaf_36_wb_clk_i _02079_ _00680_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11527_ net2069 net487 _06782_ net503 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09917__A _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14246_ clknet_leaf_75_wb_clk_i _02010_ _00611_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08007__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\] vssd1
+ vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11458_ net649 _06583_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11658__S net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] _06140_ vssd1 vssd1
+ vccd1 vccd1 _06233_ sky130_fd_sc_hd__nor2_1
XANTENNA__08102__S1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14177_ clknet_leaf_1_wb_clk_i _01941_ _00542_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ net715 net268 net697 vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11562__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ net1351 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13059_ net1267 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
Xhold1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\] vssd1
+ vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout1360 net1363 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__buf_4
Xfanout1371 net1372 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__buf_4
Xfanout1382 net1383 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__buf_4
Xfanout1393 net1394 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__buf_4
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ net815 _03560_ _03561_ _03553_ _03556_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07551_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\] net777
+ net748 _03492_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a211o_1
XANTENNA__11617__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07482_ net1139 _03419_ _03421_ _03423_ net717 vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__a41o_1
XFILLER_0_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09221_ _03641_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13936__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ net437 net429 _04444_ net544 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__o31a_1
XANTENNA__08246__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08103_ net1153 _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11250__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09083_ net1056 _05022_ _05023_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09181__A2_N _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08034_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\]
+ net894 _03975_ net1146 vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__o311a_1
Xinput70 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09827__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput81 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_1
Xhold810 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\] vssd1
+ vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold821 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\] vssd1
+ vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10980__B net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput92 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
Xhold832 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\] vssd1
+ vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07206__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13349__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold843 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\] vssd1
+ vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold854 team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\] vssd1
+ vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1124_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\] vssd1
+ vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\] vssd1
+ vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09038__S net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold887 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\] vssd1
+ vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11553__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold898 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\] vssd1
+ vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _05870_ net1670 net287 vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08936_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[971\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\] net1059
+ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__a221o_1
XANTENNA__10108__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _02937_ net559 net549 vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__and3_1
XANTENNA__11019__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\]
+ net885 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08798_ net442 net434 _04739_ net549 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o31a_1
XANTENNA__14711__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07749_ net739 _03689_ _03690_ net802 vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ _05784_ net602 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__nand2_1
XANTENNA__11035__C net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ _04820_ _05341_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10691_ net604 _06318_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10647__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11332__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08625__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ net1336 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12033__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11051__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08332__S1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ net1247 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11792__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ clknet_leaf_90_wb_clk_i _01864_ _00465_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\]
+ sky130_fd_sc_hd__dfrtp_1
X_11312_ _06469_ net2857 net409 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__mux2_1
X_15080_ net1461 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__09737__A _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12292_ net1311 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14031_ clknet_leaf_102_wb_clk_i _01795_ _00396_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ net303 net713 net825 vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07257__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net497 net647 _06666_ net417 net1877 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _04532_ net671 vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06971__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14933_ clknet_leaf_123_wb_clk_i _02688_ _01298_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10056_ net31 net1032 net906 net2843 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__o22a_1
XANTENNA__09903__C _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08173__B1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14864_ clknet_leaf_55_wb_clk_i net2346 _01229_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07920__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13815_ clknet_leaf_74_wb_clk_i _01579_ _00180_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\]
+ sky130_fd_sc_hd__dfrtp_1
X_14795_ clknet_leaf_62_wb_clk_i _02559_ _01160_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10807__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13746_ clknet_leaf_101_wb_clk_i _01510_ _00111_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10958_ net684 _05784_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08816__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09411__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11480__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13677_ clknet_leaf_105_wb_clk_i _01441_ _00042_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10889_ _06483_ net2392 net523 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12628_ net1320 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
XANTENNA__12024__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11232__A0 _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12559_ net1388 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10586__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold106 _02612_ vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\] vssd1
+ vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\] vssd1
+ vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13169__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\] vssd1
+ vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14229_ clknet_leaf_71_wb_clk_i _01993_ _00594_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07739__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08936__C1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08400__A1 net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_4
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout619 net626 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ net585 _05710_ _05711_ net359 vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o22a_1
X_06982_ _02807_ _02811_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__nor2_1
XANTENNA__10024__C _05898_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ _04657_ _04662_ net869 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11838__A2 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_2
X_08652_ _04566_ _04593_ net557 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10510__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__B1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07603_ net1158 _03543_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08583_ net1199 _04521_ _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11851__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07534_ _03473_ _03475_ net803 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06945__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__S0 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08467__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__S net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07465_ _03405_ _03406_ net812 vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout332_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1074_A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ net529 _03491_ _05144_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__nand3_2
XFILLER_0_107_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12015__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07396_ _03336_ _03337_ net743 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__mux2_1
XANTENNA__11223__A0 _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ net585 _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10991__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1241_A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10577__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1339_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ net1215 _05006_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\] net788
+ net751 _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\] vssd1
+ vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 team_03_WB.instance_to_wrap.core.register_file.registers_state\[548\] vssd1
+ vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold662 team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\] vssd1
+ vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08927__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\] vssd1
+ vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 team_03_WB.instance_to_wrap.core.register_file.registers_state\[921\] vssd1
+ vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold695 team_03_WB.instance_to_wrap.core.register_file.registers_state\[553\] vssd1
+ vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _05888_ net1708 net292 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
X_08919_ net844 _04847_ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07805__A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09899_ net359 _05735_ _05839_ _05840_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a211oi_1
XANTENNA__11829__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15172__1553 vssd1 vssd1 vccd1 vccd1 _15172__1553/HI net1553 sky130_fd_sc_hd__conb_1
XANTENNA__11181__C_N net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11930_ _06627_ net2647 net373 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10231__A _03864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ net299 net2401 net384 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__mux2_1
XANTENNA__11046__B net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13600_ net1274 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
X_10812_ net279 net2750 net521 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14580_ clknet_leaf_93_wb_clk_i _02344_ _00945_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08458__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11792_ net2231 _06622_ net334 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XANTENNA__10885__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ net1279 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XANTENNA__07540__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10743_ net1608 net531 net526 _06363_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07666__C1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07130__A1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13462_ net1395 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
X_10674_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] team_03_WB.instance_to_wrap.core.pc.current_pc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__o211a_1
XANTENNA_input95_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ net910 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_1
X_12413_ net1381 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07418__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ net1308 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10568__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11765__A1 net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15132_ net1513 vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XANTENNA__09467__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ net1368 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07433__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15063_ net1444 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ net1259 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14757__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ clknet_leaf_58_wb_clk_i _01778_ _00379_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08918__C1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11226_ net296 net2448 net492 vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08394__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11157_ net705 net272 net699 vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07715__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _04770_ net659 _05951_ _03060_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a211o_1
X_11088_ net827 net273 vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__and2_1
XANTENNA__11237__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ net18 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1
+ vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
X_14916_ clknet_leaf_125_wb_clk_i _02671_ _01281_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08697__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09894__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14847_ clknet_leaf_54_wb_clk_i net2071 _01212_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11671__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14778_ clknet_leaf_62_wb_clk_i _02542_ _01143_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13729_ clknet_leaf_0_wb_clk_i _01493_ _00094_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07250_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\] net774
+ net730 _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11205__A0 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07181_ net1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\]
+ net754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\] net724
+ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11122__D net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11756__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08621__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10964__C1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08909__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout405 _06718_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_8
Xfanout416 _06684_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout427 net428 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_8
XANTENNA__11846__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09822_ _04777_ _05762_ _05763_ _05761_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__a31o_1
Xfanout438 _04075_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12531__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout449 _06816_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__buf_4
XANTENNA__10731__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ net1018 _03724_ _04820_ _05692_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__a221o_1
X_06965_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\] net1146
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _04632_ _04645_ _04097_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_4
X_09684_ _03988_ _04178_ _04816_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a21o_1
XANTENNA__08232__S0 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06896_ _02794_ _02815_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__nor2_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08635_ net1214 _04574_ _04575_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and3_1
XANTENNA__11692__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__A _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11581__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1191_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1289_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ net934 _04506_ _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07517_ _03430_ _03458_ net612 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__mux2_4
XFILLER_0_92_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08497_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout714_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10798__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09986__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07448_ net1178 net1016 net682 vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08860__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07663__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07379_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11747__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ net1058 _05056_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11610__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08073__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ net305 net304 _06216_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__a211o_1
XANTENNA__07415__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08612__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09049_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\] net926
+ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a221o_1
X_12060_ _06626_ net2834 net361 vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__mux2_1
Xhold470 net127 vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07179__A1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold481 team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\] vssd1
+ vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net274 net704 net823 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__and3_1
Xhold492 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\] vssd1
+ vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10183__A0 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10660__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06926__A1 net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout950 net968 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__clkbuf_4
Xfanout961 net967 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__clkbuf_4
Xfanout972 net993 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_2
Xfanout983 net993 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ net1367 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\] vssd1
+ vssd1 vccd1 vccd1 net2754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ clknet_leaf_40_wb_clk_i _02465_ _01066_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\] vssd1
+ vssd1 vccd1 vccd1 net2765 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ _06614_ net2693 net376 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\] vssd1
+ vssd1 vccd1 vccd1 net2776 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11683__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ net1372 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14632_ clknet_leaf_34_wb_clk_i _02396_ _00997_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\]
+ sky130_fd_sc_hd__dfstp_1
X_11844_ _06409_ net2206 net381 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ clknet_leaf_25_wb_clk_i _02327_ _00928_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07701__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ _06608_ net482 net339 net2364 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10726_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] _05611_ net601 vssd1
+ vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__mux2_1
X_13514_ net1271 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14494_ clknet_leaf_58_wb_clk_i _02258_ _00859_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ net1400 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10657_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] team_03_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ net839 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
XANTENNA__09909__B _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13376_ net1422 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
X_10588_ net1815 net536 net597 _03103_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
X_12327_ net1390 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
X_15115_ net1496 vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15046_ net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09925__A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12258_ net1374 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11666__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ net274 net2534 net491 vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ net1656 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06917__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07445__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07164__B _03104_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08975__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07342__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ net857 _04358_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13182__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11426__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08351_ _04287_ _04292_ net868 vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07302_ _03208_ _03243_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\]
+ net969 vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08842__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07233_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\] net794
+ net730 _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_93_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11729__A1 _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11908__D_N net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15171__1552 vssd1 vssd1 vccd1 vccd1 _15171__1552/HI net1552 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07164_ _03066_ _03104_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__nand2_1
XANTENNA__08055__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08442__C _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07095_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\]
+ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__and2_1
XANTENNA__08070__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1037_A _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11576__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__C1 _05492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1204_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _05249_ _05250_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nand2b_1
Xfanout268 _06541_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_2
X_07997_ net745 _03937_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o21ai_1
Xfanout279 _06418_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
XANTENNA_fanout664_A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ _05662_ _05677_ net583 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__and3b_1
X_06948_ net612 _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09667_ net577 _05532_ _05602_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout831_A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06879_ _02799_ _02801_ _02810_ _02812_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XANTENNA__07333__A1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13092__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout929_A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11417__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ net1199 _04483_ _04490_ net844 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a211o_1
XANTENNA__09086__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11968__A1 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07097__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12090__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net2251 net488 _06794_ net512 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a22o_1
XANTENNA__11043__C net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11432__A3 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07192__S0 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ net2017 net1023 net1019 team_03_WB.instance_to_wrap.CPU_DAT_I\[28\] vssd1
+ vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire614 _02842_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10640__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11491_ _06612_ net2573 net393 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__mux2_1
XANTENNA__10655__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13230_ net1281 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
X_10442_ net305 net304 _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08597__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ net1248 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
X_10373_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] _06145_ vssd1 vssd1
+ vccd1 vccd1 _06204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12112_ net1135 net1739 net1997 _06282_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input58_A gpio_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ net1307 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12043_ _06612_ net2744 net361 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07265__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07572__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout780 net783 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout791 net796 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ clknet_leaf_4_wb_clk_i _01758_ _00359_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ net1305 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
XANTENNA__07324__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ net1298 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11408__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14615_ clknet_leaf_76_wb_clk_i _02379_ _00980_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__09077__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11827_ net646 _06659_ net458 net328 net2096 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a32o_1
XANTENNA__11959__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07088__B1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08824__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14546_ clknet_leaf_100_wb_clk_i _02310_ _00911_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07627__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ _06584_ net465 net339 net2509 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
XANTENNA__12081__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _05500_ _05932_ net604 vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10631__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14477_ clknet_leaf_106_wb_clk_i _02241_ _00842_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12346__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11689_ _06731_ net385 net344 net2161 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ net1308 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11187__A2 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13359_ net1283 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08052__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__S net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10934__A2 _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07260__B1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ net1141 _03857_ _03859_ _03861_ net719 vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13177__A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15029_ clknet_leaf_55_wb_clk_i _02749_ _01394_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09001__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07851_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[763\] net748
+ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__o221a_1
XANTENNA__10698__B2 _06336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07563__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_07782_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02821_ _03107_ vssd1
+ vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a21o_2
XFILLER_0_39_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09521_ _04829_ _05462_ _02993_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07315__A1 net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08512__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _05111_ _05128_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07622__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\]
+ net991 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09068__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ _05323_ _05324_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13640__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08334_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08276__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06953__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10983__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10622__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10083__C1 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ _04193_ _04206_ net845 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_8
XANTENNA_fanout412_A _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11160__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07216_ _03156_ _03157_ net737 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__mux2_1
XANTENNA__08579__B1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07147_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\] net733
+ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08043__A2 _02821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1321_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__C_N _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1419_A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07251__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ net1124 _03018_ net1157 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout781_A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14818__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10138__A0 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
Xfanout1019 net1022 vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11886__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__C net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14968__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11638__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _05239_ _05271_ _05273_ _05231_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__a31o_1
X_10991_ net1242 net827 _06414_ net666 vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07306__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11335__A _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ net1371 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12661_ net1268 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14400_ clknet_leaf_133_wb_clk_i _02164_ _00765_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\]
+ sky130_fd_sc_hd__dfrtp_1
X_11612_ _06686_ net385 net353 net2457 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12592_ net1427 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14331_ clknet_leaf_27_wb_clk_i _02095_ _00696_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ net494 net616 _06653_ net486 net1867 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a32o_1
XANTENNA__10385__S net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11810__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11070__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08019__C1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14262_ clknet_leaf_85_wb_clk_i _02026_ _00627_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11474_ net2415 net399 _06772_ net512 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
XANTENNA__07490__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11169__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ net1381 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10425_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] _06138_ vssd1 vssd1
+ vccd1 vccd1 _06246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14193_ clknet_leaf_94_wb_clk_i _01957_ _00558_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10916__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ net1369 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10356_ _06098_ _06189_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14498__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07793__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08990__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ net1266 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
X_10287_ _04475_ _02766_ net671 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12026_ _06768_ net461 net366 net2374 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__a22o_1
XANTENNA__09534__A2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07426__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08742__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__B _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07640__S1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A3 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15170__1551 vssd1 vssd1 vccd1 vccd1 _15170__1551/HI net1551 sky130_fd_sc_hd__conb_1
X_13977_ clknet_leaf_103_wb_clk_i _01741_ _00342_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11245__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12928_ net1379 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12859_ net1344 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10604__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14529_ clknet_leaf_0_wb_clk_i _02293_ _00894_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09470__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07076__A3 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08050_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\] net767
+ net742 _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13715__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07001_ _02939_ _02941_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09385__A _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07233__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08430__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08981__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ net443 net435 _04893_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nor3_1
XANTENNA__13865__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\] net749
+ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__a221o_1
XANTENNA__11868__A0 _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ net442 net434 _04807_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__or3_1
XANTENNA__07536__A1 net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07834_ net816 _03775_ net720 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10540__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A3 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07765_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\]
+ net874 _03706_ net1143 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout362_A _06818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11155__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ _03823_ _04444_ net664 _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08497__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ _03620_ _03621_ _03629_ _03637_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__o22a_4
XFILLER_0_91_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09435_ _05375_ _05376_ net558 vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__mux2_1
XANTENNA__10994__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1271_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout627_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1369_A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _05185_ _05191_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\]
+ net983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\] net1217
+ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09297_ _04619_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09994__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\]
+ net948 net1065 vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout996_A _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08179_ net551 _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10210_ _02889_ _06039_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07224__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07808__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08421__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ net654 net706 net268 net697 vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11571__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _05981_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_41_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XANTENNA__14790__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07019__S net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11859__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11049__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _02811_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nor3_1
X_13900_ clknet_leaf_5_wb_clk_i _01664_ _00265_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\]
+ sky130_fd_sc_hd__dfrtp_1
X_14880_ clknet_leaf_52_wb_clk_i _02643_ _01245_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10531__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13831_ clknet_leaf_69_wb_clk_i _01595_ _00196_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09819__A3 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13762_ clknet_leaf_130_wb_clk_i _01526_ _00127_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ net313 net311 net322 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12713_ net1250 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13693_ clknet_leaf_67_wb_clk_i _01457_ _00058_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12036__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ net1314 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ net1377 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10062__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ clknet_leaf_2_wb_clk_i _02078_ _00679_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\]
+ sky130_fd_sc_hd__dfrtp_1
X_11526_ net652 _06638_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08660__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11939__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ net494 net615 _06582_ net397 net2107 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a32o_1
X_14245_ clknet_leaf_107_wb_clk_i _02009_ _00610_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10408_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] net678 _06230_ _06232_
+ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__o22a_1
X_14176_ clknet_leaf_132_wb_clk_i _01940_ _00541_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08313__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ net510 net631 _06746_ net407 net1978 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13127_ net1399 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
X_10339_ _06112_ _06115_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10144__A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06974__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__A _03821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ net1347 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XANTENNA__11674__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1352 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__buf_4
X_12009_ _06759_ net462 net365 net2579 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a22o_1
Xfanout1361 net1363 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__buf_2
XANTENNA__10522__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1372 net1373 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__buf_4
XANTENNA__08191__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1383 net1386 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__clkbuf_2
Xfanout1394 net1406 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__buf_2
XFILLER_0_108_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\]
+ net882 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08479__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14513__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07481_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\] net789
+ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ _03280_ _03314_ _05160_ net605 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12027__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09151_ net579 _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08102_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\]
+ net764 net1119 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09082_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\]
+ net963 net1067 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__mux4_1
XANTENNA__11250__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11849__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\]
+ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold800 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\] vssd1
+ vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xinput60 gpio_in[35] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xinput71 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold811 team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\] vssd1
+ vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput93 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold822 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\] vssd1
+ vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11002__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07628__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\] vssd1
+ vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_03_WB.instance_to_wrap.ADR_I\[15\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08223__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold855 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\] vssd1
+ vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07757__A1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold866 team_03_WB.instance_to_wrap.core.register_file.registers_state\[833\] vssd1
+ vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11553__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold877 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\] vssd1
+ vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 net130 vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _05869_ net1831 net287 vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__mux2_1
Xhold899 team_03_WB.instance_to_wrap.core.register_file.registers_state\[901\] vssd1
+ vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1117_A _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ _04875_ _04876_ net864 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10989__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10513__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ net549 _04807_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08182__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08459__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07817_ _03756_ _03758_ net609 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__mux2_1
X_08797_ net843 _04738_ _04727_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_93_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07390__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09989__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14193__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07748_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\]
+ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08893__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ net816 _03614_ net717 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12709__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _04268_ _04355_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] _06317_ vssd1 vssd1
+ vccd1 vccd1 _06330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07693__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ _05285_ _05290_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_105_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ net1285 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
XANTENNA__11051__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07996__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ _06454_ net2649 net409 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XANTENNA__09737__B _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12291_ net1300 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XANTENNA__12444__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14030_ clknet_leaf_72_wb_clk_i _01794_ _00395_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11242_ net496 net617 _06688_ net413 net2303 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11173_ net1038 net831 net270 net666 vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06956__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] net671 vssd1 vssd1 vccd1
+ vccd1 _05966_ sky130_fd_sc_hd__nand2_1
XANTENNA_input40_A gpio_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11494__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14932_ clknet_leaf_125_wb_clk_i _02687_ _01297_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10055_ net32 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1
+ vccd1 vccd1 _02676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08173__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ clknet_leaf_54_wb_clk_i net1652 _01228_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07920__A1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13814_ clknet_leaf_84_wb_clk_i _01578_ _00179_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14794_ clknet_leaf_61_wb_clk_i _02558_ _01159_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ clknet_leaf_96_wb_clk_i _01509_ _00110_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[3\] net308 net684 vssd1
+ vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12009__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07684__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13676_ clknet_leaf_9_wb_clk_i _01440_ _00041_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10888_ _06480_ _06481_ _06482_ net586 vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__o211a_4
XFILLER_0_94_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12627_ net1260 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
XANTENNA__08859__S0 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07436__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10035__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12558_ net1340 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XANTENNA__08633__C1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11669__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ _06505_ net2796 net395 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold107 team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\] vssd1
+ vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12489_ net1247 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold118 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\] vssd1
+ vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11941__D_N net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\] vssd1
+ vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14228_ clknet_leaf_95_wb_clk_i _01992_ _00593_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08936__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159_ clknet_leaf_99_wb_clk_i _01923_ _00524_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout609 _02843_ vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09663__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06981_ net612 _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a21oi_2
XANTENNA__13185__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ net1061 _04660_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08279__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
X_08651_ net441 net433 _04592_ net548 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__o31a_1
Xfanout1191 net1196 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07911__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ net1127 _03539_ _03540_ _03542_ net1113 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__a311o_1
XFILLER_0_90_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08582_ net934 _04523_ _04522_ net1057 vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__o211a_1
XANTENNA__11136__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07533_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\] net775
+ net750 _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08011__S1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07464_ net1108 _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ net529 _03491_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__and3_1
XANTENNA__11152__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07395_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\]
+ net769 vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ net529 _02948_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__and3_1
XANTENNA__09838__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10991__B net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07522__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11774__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09065_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\] net926
+ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1234_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08016_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[689\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\] vssd1
+ vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold641 team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\] vssd1
+ vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout694_A _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08927__B1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\] vssd1
+ vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 team_03_WB.instance_to_wrap.ADR_I\[21\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold674 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\] vssd1
+ vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1401_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\] vssd1
+ vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold696 team_03_WB.instance_to_wrap.core.register_file.registers_state\[410\] vssd1
+ vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07792__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ _03788_ net660 vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout861_A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net866 _04859_ _04854_ net846 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__o211a_1
X_09898_ net325 _05397_ _05403_ _05513_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ net1063 _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07902__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11860_ net271 net2278 net381 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09104__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _06415_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10658__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ net2204 _06479_ net335 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09655__A1 _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11343__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13530_ net1278 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
XANTENNA__07666__B1 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] _05686_ net603 vssd1
+ vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11462__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13461_ net1333 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
X_10673_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ net911 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07418__B1 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ net1350 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08615__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ net1308 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
XANTENNA_input88_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11489__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15131_ net1512 vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
X_12343_ net1417 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XANTENNA__07268__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15062_ net1443 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
X_12274_ net1410 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14013_ clknet_leaf_66_wb_clk_i _01777_ _00378_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11225_ net2632 net492 _06683_ net512 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
XANTENNA__10725__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08394__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ net2119 net417 _06655_ net500 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a22o_1
XANTENNA__06900__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] net659 vssd1 vssd1 vccd1
+ vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11087_ _06469_ net2419 net421 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14915_ clknet_leaf_125_wb_clk_i _02670_ _01280_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10038_ net19 net1033 net907 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1
+ vccd1 vccd1 _02693_ sky130_fd_sc_hd__o22a_1
XANTENNA__11237__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ clknet_leaf_55_wb_clk_i _02610_ _01211_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14777_ clknet_leaf_61_wb_clk_i _02541_ _01142_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11989_ _06753_ net465 net449 net2397 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11253__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13728_ clknet_leaf_133_wb_clk_i _01492_ _00093_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11453__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07121__A2 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13659_ clknet_leaf_28_wb_clk_i _01423_ _00024_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07409__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07180_ _03116_ _03121_ net816 vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08562__A _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11399__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08082__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07424__A3 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07178__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08909__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout406 _06718_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout417 _06635_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_6
XFILLER_0_61_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09821_ net572 _05114_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__or2_1
XANTENNA__08501__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 _06560_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_8
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_2
XANTENNA__07593__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09752_ _03727_ net588 _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a21oi_1
X_06964_ _02900_ _02905_ net818 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__mux2_1
X_08703_ _04639_ _04644_ net869 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__mux2_1
X_09683_ _05298_ _05597_ _05296_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__a21o_1
X_06895_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] net1015 _02836_
+ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or3_4
XANTENNA__08232__S1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__S net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_A _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10495__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07896__B1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\]
+ net979 net1072 vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10986__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09098__C1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[189\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\] net967 net918
+ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12259__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1184_A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ net719 _03441_ _03450_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__o22a_4
XFILLER_0_119_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08496_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\]
+ net989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\] net1075
+ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__o221a_1
XANTENNA__11444__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07112__A2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07447_ net720 _03382_ _03388_ _03373_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o31a_4
XANTENNA__10798__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1351_A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07378_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\] net729
+ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11747__A2 _06569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ net1209 _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and3_1
XANTENNA__11610__B net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08073__B1 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\] net942
+ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13949__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold460 team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\] vssd1
+ vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold471 _02634_ vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ net2533 net425 _06578_ net501 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a22o_1
Xhold482 team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\] vssd1
+ vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\] vssd1
+ vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net945 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout951 net953 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
Xfanout962 net964 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout984 net987 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout995 net996 vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_4
XANTENNA__11057__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ net1268 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
XANTENNA__09876__A1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\] vssd1
+ vssd1 vccd1 vccd1 net2744 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ clknet_leaf_40_wb_clk_i _02464_ _01065_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\] vssd1
+ vssd1 vccd1 vccd1 net2755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\] vssd1
+ vssd1 vccd1 vccd1 net2766 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _06613_ net2815 net373 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
XANTENNA__09750__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\] vssd1
+ vssd1 vccd1 vccd1 net2777 sky130_fd_sc_hd__dlygate4sd3_1
X_12892_ net1340 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ clknet_leaf_63_wb_clk_i _02395_ _00996_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_115_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09089__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net281 net2128 net382 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ clknet_leaf_129_wb_clk_i _02326_ _00927_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ _06607_ net478 net338 net2307 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a22o_1
XANTENNA__08300__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13513_ net1325 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10725_ net525 _06353_ _06354_ net533 net2031 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a32o_1
XFILLER_0_138_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14493_ clknet_leaf_66_wb_clk_i _02257_ _00858_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13444_ net1395 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__A _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11199__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\] team_03_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ net839 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11738__A2 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13375_ net1402 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
X_10587_ net1829 net536 net597 _03059_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10946__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ net1495 vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_2
X_12326_ net1419 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
XANTENNA__07811__B1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14874__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15045_ net171 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09159__A3 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09925__B _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ net1288 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__inv_2
X_11208_ _06442_ net2411 net491 vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__mux2_1
X_12188_ net1636 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10152__A _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ net2254 net420 _06645_ net515 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08119__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09941__A _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09867__B2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07878__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14829_ clknet_leaf_40_wb_clk_i net1807 _01194_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09619__B2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07893__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08350_ net1210 _04290_ _04291_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ _03241_ _03242_ _02843_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08281_ _04217_ _04222_ net870 vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07232_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08055__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07163_ _03066_ _03104_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__and2_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _03027_ _03030_ _03035_ net1110 net1131 vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__o221a_1
XANTENNA__07802__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_62_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09004__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08358__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07636__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07566__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11362__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _02954_ _05735_ _05745_ _05733_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__a211oi_4
XANTENNA__07030__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout269 _06532_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\]
+ net798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[688\] net735
+ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07581__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__A net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ _05227_ _05660_ _05217_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__a21o_1
XANTENNA__11114__A0 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06947_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] _02808_ _02818_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout657_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1399_A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ _05513_ _05521_ _05522_ net325 _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a221o_1
X_06878_ _02800_ _02802_ _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__o22a_4
X_08617_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ _05371_ _05523_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout824_A _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09997__S net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10001__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _04486_ _04489_ net1199 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07097__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08479_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\]
+ net988 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\] net926
+ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__o221a_1
XFILLER_0_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10510_ net157 net1023 net1019 net1987 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
X_15139__1520 vssd1 vssd1 vccd1 vccd1 _15139__1520/HI net1520 sky130_fd_sc_hd__conb_1
XANTENNA__07192__S1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11490_ _06611_ net2756 net393 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14897__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ _06028_ _06056_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08597__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10372_ net286 _06089_ _06202_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13160_ net1351 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08061__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ net1135 net1687 net2086 _06302_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13091_ net1262 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09546__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12042_ _06611_ net2866 net361 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__mux2_1
Xhold290 _02583_ vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10156__A1 _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11068__A net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout770 net772 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_2
Xfanout781 net783 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14277__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout792 net793 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07309__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13993_ clknet_leaf_60_wb_clk_i _01757_ _00358_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09849__A1 _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ net1416 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11656__A1 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08521__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08521__B2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12875_ net1254 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
X_14614_ clknet_leaf_85_wb_clk_i _02378_ _00979_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\]
+ sky130_fd_sc_hd__dfstp_1
X_11826_ _06658_ net481 net330 net2393 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11234__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09904__C_N _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07088__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ clknet_leaf_93_wb_clk_i _02309_ _00910_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11757_ net646 _06582_ net457 net337 net2093 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10708_ _06149_ net600 _06315_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14476_ clknet_leaf_8_wb_clk_i _02240_ _00841_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _06730_ net385 net344 net1955 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13427_ net1309 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10639_ net1145 net2879 net839 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XANTENNA__10919__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13358_ net1279 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XANTENNA__10395__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__A0 _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13458__A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12309_ net1267 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XANTENNA__07260__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13289_ net1332 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15028_ clknet_leaf_56_wb_clk_i _02748_ _01393_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07456__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11344__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07850_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__or3_1
XANTENNA__11895__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07781_ _03700_ _03701_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__o21a_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_09520_ net568 _05459_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13193__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ _05391_ _05392_ net558 vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07720__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08402_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\] net927
+ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__a221o_1
X_09382_ _04354_ _05322_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08333_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08276__B1 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07079__B2 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08264_ net863 _04204_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11160__B _06657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07215_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\]
+ net753 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__mux2_1
X_08195_ _04135_ _04136_ net855 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout405_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1147_A team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07146_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\]
+ net879 _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09846__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11583__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11587__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07077_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[386\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\]
+ net772 net1129 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1314_A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07539__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11886__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07979_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\] net798
+ _02869_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout941_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _05239_ _05271_ _05273_ _05232_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a31o_1
X_10990_ net2713 net425 _06566_ net496 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XANTENNA__07937__S0 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__C1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09649_ _03428_ _04295_ net664 _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07711__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12660_ net1320 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11611_ _06685_ net388 net355 net2496 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XANTENNA__08267__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ net1389 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11351__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ clknet_leaf_20_wb_clk_i _02094_ _00695_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ net494 net616 _06652_ net486 net2092 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11070__B net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07490__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14261_ clknet_leaf_71_wb_clk_i _02025_ _00626_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11473_ net655 _06598_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input70_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net1352 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
X_10424_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _06245_ net678 vssd1
+ vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ clknet_leaf_113_wb_clk_i _01956_ _00557_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08034__A3 net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__C1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10916__A3 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ net1411 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10355_ _06100_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08990__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13074_ net1420 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
X_10286_ _05971_ _05973_ _06126_ _05968_ _05965_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a311o_1
XANTENNA__11326__A0 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12025_ net627 _06588_ net465 net366 net2314 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__a32o_1
XANTENNA__11877__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__C _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ clknet_leaf_10_wb_clk_i _01740_ _00341_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11245__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12927_ net1375 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10852__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ net1371 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
XANTENNA__08835__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11809_ _06634_ _06803_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__or2_1
XANTENNA__12357__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12789_ net1267 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14528_ clknet_leaf_134_wb_clk_i _02292_ _00893_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14459_ clknet_leaf_35_wb_clk_i _02223_ _00824_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] _02928_ net683 _02941_
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10368__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11565__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14442__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07769__C1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08430__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11200__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08951_ net843 _04871_ _04877_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__a31o_4
XANTENNA__11317__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07902_ net815 _03833_ _03843_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08882_ _04080_ _04807_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08733__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09605__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _03773_ _03774_ net1107 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11436__A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\]
+ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ net541 _05443_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07695_ net1138 _03632_ _03634_ _03636_ net717 vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__a41o_1
XANTENNA__11870__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ net547 _04894_ _04955_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_71_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06964__S net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10994__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _05193_ _05305_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11171__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08316_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[920\] net1009
+ _04252_ net1064 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09296_ _03459_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07472__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\]
+ net946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1431_A net1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__B2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08178_ net439 net430 _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout891_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout989_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08421__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\]
+ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10140_ _03390_ _05980_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08972__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_101_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10071_ team_03_WB.instance_to_wrap.core.i_hit _05914_ vssd1 vssd1 vccd1 vccd1 _05915_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_41_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11049__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13830_ clknet_leaf_74_wb_clk_i _01594_ _00195_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ clknet_leaf_0_wb_clk_i _01525_ _00126_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10973_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\] net315 net310 net319
+ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__or4_1
XANTENNA__11780__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__A_N net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13561__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12712_ net1351 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13692_ clknet_leaf_119_wb_clk_i _01456_ _00057_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_108_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ net1300 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12574_ net1385 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07999__C1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14313_ clknet_leaf_49_wb_clk_i _02077_ _00678_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11525_ net2238 net486 _06781_ net496 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XANTENNA__08660__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14244_ clknet_leaf_20_wb_clk_i _02008_ _00609_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\]
+ sky130_fd_sc_hd__dfrtp_1
X_11456_ net495 net615 _06581_ net397 net2243 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08007__A3 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10407_ net285 _06231_ net678 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ clknet_leaf_117_wb_clk_i _01939_ _00540_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\]
+ sky130_fd_sc_hd__dfrtp_1
X_11387_ net1243 net834 _06536_ net667 vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ net1426 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
X_10338_ _06150_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06974__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09933__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ net1287 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
X_10269_ _06107_ _06109_ _05976_ _05979_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__a211o_1
XANTENNA__08176__C1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1340 net1342 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__buf_4
XFILLER_0_108_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12008_ _06758_ net471 net368 net2536 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a22o_1
Xfanout1351 net1352 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__buf_4
Xfanout1362 net1363 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__buf_4
Xfanout1373 net1387 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__buf_2
Xfanout1384 net1385 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__buf_4
Xfanout1395 net1396 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__buf_4
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10160__A _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13959_ clknet_leaf_66_wb_clk_i _01723_ _00324_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08479__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07480_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\] net762
+ net1011 vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21a_1
XANTENNA__10825__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09979__A0 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10038__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _05084_ _05086_ _05089_ _05091_ net556 net566 vssd1 vssd1 vccd1 vccd1 _05092_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08100__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[474\]
+ net765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\] net1143
+ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07454__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[461\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\] net1202
+ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__o221a_1
XANTENNA__11250__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08032_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\]
+ net894 _03973_ net1122 vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__o311a_1
Xinput50 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 gpio_in[5] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
Xinput72 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold801 team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\] vssd1
+ vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold812 team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\] vssd1
+ vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold823 team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\] vssd1
+ vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07206__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput83 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_1
Xinput94 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11002__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold834 team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\] vssd1
+ vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\] vssd1
+ vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_03_WB.instance_to_wrap.core.register_file.registers_state\[497\] vssd1
+ vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\] vssd1
+ vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\] vssd1
+ vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09983_ _05868_ net1915 net287 vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__mux2_1
Xhold889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\] vssd1
+ vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ net1213 _04872_ _04873_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout1012_A _02821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__C1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ net844 _04787_ _04793_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ net1178 _02814_ _02924_ net1246 _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_135_1403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08796_ _04730_ _04731_ _04737_ _04734_ net1059 _02788_ vssd1 vssd1 vccd1 vccd1 _04738_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__08178__C _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07747_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout737_A net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10816__A2 _06420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08475__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _03618_ _03619_ net812 vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14488__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ _03064_ _05357_ _05358_ net571 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__o211a_1
XANTENNA__12018__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout904_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11105__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ _05288_ _05289_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__and2_1
XANTENNA__11332__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09279_ _04893_ _05219_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__xor2_1
XFILLER_0_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08922__B net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ _06620_ net2819 net409 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08414__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ net1353 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ net1241 net831 net279 net668 vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11172_ net2157 net419 _06665_ net506 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
XANTENNA__06956__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__inv_2
XANTENNA__12460__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14931_ clknet_leaf_126_wb_clk_i _02686_ _01296_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10054_ net33 net1032 net906 net2850 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__o22a_1
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__A1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ clknet_leaf_54_wb_clk_i net1788 _01227_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09502__A1_N team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13813_ clknet_leaf_89_wb_clk_i _01577_ _00178_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13705__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14793_ clknet_leaf_40_wb_clk_i _02557_ _01158_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13744_ clknet_leaf_81_wb_clk_i _01508_ _00109_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10956_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[3\] net306 vssd1 vssd1
+ vccd1 vccd1 _06538_ sky130_fd_sc_hd__and2_1
XANTENNA__07133__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13675_ clknet_leaf_45_wb_clk_i _01439_ _00040_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11480__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ net685 _05811_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12626_ net1420 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08859__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11768__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12557_ net1318 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XANTENNA__08633__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _06626_ net2641 net393 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12488_ net1285 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[3\] vssd1 vssd1 vccd1
+ vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold119 team_03_WB.instance_to_wrap.CPU_DAT_I\[2\] vssd1 vssd1 vccd1 vccd1 net1703
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ clknet_leaf_108_wb_clk_i _01991_ _00592_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ net2468 net397 _06759_ net501 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08936__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14158_ clknet_leaf_70_wb_clk_i _01922_ _00523_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07295__S0 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13109_ net1262 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
X_14089_ clknet_leaf_59_wb_clk_i _01853_ _00454_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\]
+ sky130_fd_sc_hd__dfrtp_1
X_06980_ net612 _02893_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07464__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1170 net1172 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1181 net1197 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07183__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08650_ _04591_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__inv_2
Xfanout1192 net1196 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07372__A0 _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07601_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[409\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\]
+ net782 net1126 vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08581_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XANTENNA__11136__D net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07532_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\]
+ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08295__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09664__A2 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ net1153 _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08872__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098__1479 vssd1 vssd1 vccd1 vccd1 _15098__1479/HI net1479 sky130_fd_sc_hd__conb_1
XFILLER_0_130_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09202_ net584 net579 net572 _05124_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__and4_2
XFILLER_0_85_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11152__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07394_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\]
+ net769 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__mux2_1
XANTENNA__11759__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _02804_ _02944_ net591 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07522__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09064_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\] net942
+ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08015_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[529\]
+ net785 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold620 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\] vssd1
+ vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10065__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold631 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\] vssd1
+ vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 net175 vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1227_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold653 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\] vssd1
+ vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold664 team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\] vssd1
+ vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\] vssd1
+ vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11595__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold686 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\] vssd1
+ vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold697 team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\] vssd1
+ vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _05887_ net1883 net293 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14160__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07374__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _04855_ _04856_ _04858_ _04857_ net935 net857 vssd1 vssd1 vccd1 vccd1 _04859_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11608__B net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ net326 _05419_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout854_A _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\]
+ net987 net1074 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07363__B1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10810_ net692 _05583_ net587 vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13878__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11790_ net2572 _06621_ net332 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux2_1
XANTENNA__07115__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__A2 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11998__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ net1881 net531 net526 _06362_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11343__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07666__A1 net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11462__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07130__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13460_ net1393 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
X_10672_ _05429_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__nand2_1
XANTENNA__08933__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12411_ net1362 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11214__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ net1309 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XANTENNA__08615__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__C1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15130_ net1511 vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12342_ net1343 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11765__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07549__A _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15061_ net1442 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
X_12273_ net1304 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__inv_2
XANTENNA__08918__A1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ clknet_leaf_120_wb_clk_i _01776_ _00377_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11224_ _06456_ _06517_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__nor2_1
XANTENNA__10725__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11155_ net628 _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ _02834_ _05916_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__or2_4
XANTENNA__07715__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ _06454_ net2405 net421 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10489__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ net20 net1036 net909 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1
+ vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
X_14914_ clknet_leaf_125_wb_clk_i _02669_ _01279_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11237__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07354__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__A2 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08551__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14845_ clknet_leaf_55_wb_clk_i net1921 _01210_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08529__S0 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__A _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14776_ clknet_leaf_40_wb_clk_i _02540_ _01141_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11988_ net273 net2667 net448 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__mux2_1
XANTENNA__11989__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11253__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07657__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ clknet_leaf_121_wb_clk_i _01491_ _00092_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08854__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[6\] net306 vssd1 vssd1
+ vccd1 vccd1 _06524_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11453__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09939__A _03526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13658_ clknet_leaf_22_wb_clk_i _01422_ _00023_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14033__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12609_ net1287 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ net1336 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11756__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08909__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09031__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout407 _06718_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_8
X_09820_ net567 _05134_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__or2_1
Xfanout418 _06635_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_4
Xfanout429 net430 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_2
XANTENNA__07593__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _04816_ _05692_ net664 vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__o21a_1
X_06963_ net1111 _02903_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a21o_1
X_08702_ net1214 _04642_ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__o21a_1
X_09682_ _05296_ _05298_ _05597_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__nand3_1
X_06894_ _02823_ _02831_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08542__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08633_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\] net1076
+ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a221o_1
XANTENNA__11692__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08564_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[29\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07515_ net820 _03456_ net723 vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11444__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ net861 _04433_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08845__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1177_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10652__A0 net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07446_ _03386_ _03387_ net812 vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout602_A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07377_ net743 _03315_ _03316_ _03317_ _03318_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09116_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\] net1203
+ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11747__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08073__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09047_ _04987_ _04988_ net852 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07281__C1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07259__S0 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\] vssd1
+ vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 team_03_WB.instance_to_wrap.core.register_file.registers_state\[282\] vssd1
+ vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\] vssd1
+ vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09573__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\] vssd1
+ vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 team_03_WB.instance_to_wrap.core.register_file.registers_state\[249\] vssd1
+ vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11380__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_2
Xfanout941 net943 vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
XANTENNA__06926__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _03136_ net660 vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__nor2_1
Xfanout952 net953 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__clkbuf_4
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
Xfanout974 net993 vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__clkbuf_4
Xfanout985 net987 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ net1409 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout996 _04085_ vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__C _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08928__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1150 team_03_WB.instance_to_wrap.core.register_file.registers_state\[118\] vssd1
+ vssd1 vccd1 vccd1 net2734 sky130_fd_sc_hd__dlygate4sd3_1
X_11911_ _06612_ net2726 net373 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__mux2_1
Xhold1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\] vssd1
+ vssd1 vccd1 vccd1 net2745 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\] vssd1
+ vssd1 vccd1 vccd1 net2756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11683__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ net1348 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
Xhold1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\] vssd1
+ vssd1 vccd1 vccd1 net2767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\] vssd1
+ vssd1 vccd1 vccd1 net2778 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ clknet_leaf_78_wb_clk_i _02394_ _00995_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10891__B1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11842_ _06455_ net465 vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09089__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ clknet_leaf_130_wb_clk_i _02325_ _00926_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07639__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11773_ net656 _06606_ net473 net339 net2129 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10643__A0 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ net1327 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
X_10724_ _05833_ net601 vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
X_14492_ clknet_leaf_126_wb_clk_i _02256_ _00857_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08663__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ net1400 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10655_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ net839 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08064__A1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11738__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13374_ net1400 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
X_10586_ net1703 net535 net596 _03023_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15113_ net1494 vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_2
XFILLER_0_23_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12325_ net1288 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
XANTENNA__07811__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15044_ clknet_leaf_56_wb_clk_i _02764_ _01409_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09494__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ net1413 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
XANTENNA__06911__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _06438_ net2385 net490 vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__mux2_1
X_12187_ net1667 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15097__1478 vssd1 vssd1 vccd1 vccd1 _15097__1478/HI net1478 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ net275 net656 net708 net699 vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09941__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _06612_ net2429 net421 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07327__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08524__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11123__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07742__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14828_ clknet_leaf_32_wb_clk_i net1859 _01193_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08827__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14759_ clknet_leaf_118_wb_clk_i _02523_ _01124_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10634__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07300_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] net821 vssd1 vssd1 vccd1
+ vccd1 _03242_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08280_ net1059 _04218_ _04219_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07231_ net1184 net877 team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\]
+ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11203__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07162_ _03075_ _03081_ _03102_ _02843_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a211o_2
XANTENNA__08055__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07093_ _03032_ _03034_ net746 vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09004__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07566__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ net327 _05403_ _05737_ _05740_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11901__A3 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\]
+ net784 vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout385_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ net583 _05663_ _05664_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a31o_4
X_06946_ _02862_ _02876_ _02887_ net718 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__o22a_4
XFILLER_0_39_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09665_ _02804_ _03139_ net539 _05604_ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_59_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout552_A _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _02808_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout1294_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08616_ net859 _04556_ _04557_ _04555_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09596_ _04778_ _05527_ _05531_ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08547_ net917 _04487_ _04488_ net1210 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout817_A _02846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11968__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ net942 _04418_ _04419_ net853 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__o211a_1
XANTENNA__12090__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13916__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07429_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\] net787
+ net1037 _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10440_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] net679 _06256_ _06258_
+ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10928__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ _05983_ _05986_ _06088_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ net1135 _06305_ _06821_ net842 vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07827__A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13090_ net1349 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09546__A1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _06609_ net2752 net364 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_1
XANTENNA__11349__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\] vssd1
+ vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\] vssd1
+ vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10156__A2 net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11783__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net785 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_4
XANTENNA__13564__A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout771 net772 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
Xfanout782 net783 vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13992_ clknet_leaf_35_wb_clk_i _01756_ _00357_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout793 net795 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07562__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12943_ net1407 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11084__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12874_ net1248 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11825_ net658 _06656_ net472 net330 net1924 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14613_ clknet_leaf_71_wb_clk_i _02377_ _00978_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11234__D net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11959__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14544_ clknet_leaf_82_wb_clk_i _02308_ _00909_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\]
+ sky130_fd_sc_hd__dfrtp_1
X_11756_ net646 _06581_ net457 net337 net2222 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a32o_1
XANTENNA__09482__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06906__A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12081__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ net2469 net531 net526 _06343_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
X_14475_ clknet_leaf_37_wb_clk_i _02239_ _00840_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11687_ _06729_ net386 net345 net2248 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13426_ net1331 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10638_ net1138 net2047 net839 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10919__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09785__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ net1318 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
X_10569_ net2005 net534 net595 _05879_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10395__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ net1322 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XANTENNA__14991__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ net1331 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15027_ clknet_leaf_41_wb_clk_i _02747_ _01392_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09537__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11259__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12239_ net1748 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11344__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07780_ _03715_ _03721_ _02864_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ _05116_ _05118_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08401_ _04341_ _04342_ net1215 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13939__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09381_ _04354_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10607__A0 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _04270_ _04271_ _04272_ _04273_ net857 net918 vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08276__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08507__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10083__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11280__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ net867 _04196_ _04199_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07214_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\]
+ net753 vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\]
+ net947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\] net929
+ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11868__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07145_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\]
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__and2_1
XANTENNA__07236__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout300_A _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1042_A net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07787__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08984__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07076_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\]
+ net878 _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1307_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07539__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08736__C1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09862__A _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout767_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__or3_1
XFILLER_0_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14714__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ _05648_ _05649_ _05657_ _05658_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__o211ai_4
X_06929_ net1145 net1152 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__nor2_8
XANTENNA__11638__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11108__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09700__A1 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10012__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net542 _05588_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__nand2_1
XANTENNA__07937__S1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09579_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11610_ net1038 net701 _06803_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__or3_1
XFILLER_0_132_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12590_ net1340 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07475__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15096__1477 vssd1 vssd1 vccd1 vccd1 _15096__1477/HI net1477 sky130_fd_sc_hd__conb_1
XANTENNA__11351__B net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net495 net619 _06651_ net486 net1855 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11810__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14260_ clknet_leaf_95_wb_clk_i _02024_ _00625_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08019__A1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ net2635 net399 _06771_ net516 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ net1360 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XANTENNA__11778__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _06242_ _06244_ net285 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__mux2_1
XANTENNA__11023__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14191_ clknet_leaf_99_wb_clk_i _01955_ _00556_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07557__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ net1345 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
X_10354_ _06101_ _06187_ _06092_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__and3b_1
XFILLER_0_81_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input63_A gpio_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13073_ net1316 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10285_ _05973_ _06126_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08727__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ _06767_ net483 net367 net2565 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__a22o_1
XANTENNA__09772__A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11629__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ clknet_leaf_74_wb_clk_i _01739_ _00340_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10837__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11245__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ net1385 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ net1357 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12638__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__B _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ net2530 _06633_ net334 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ net1322 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11261__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09012__A _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11739_ net2122 net268 net342 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
X_14527_ clknet_leaf_114_wb_clk_i _02291_ _00892_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09947__A _03389_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07481__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ clknet_leaf_8_wb_clk_i _02222_ _00823_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09758__A1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ net1422 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XANTENNA__09758__B2 _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14389_ clknet_leaf_89_wb_clk_i _02153_ _00754_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10368__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11565__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07233__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08950_ net847 _04884_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08997__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ net819 _03838_ _03840_ _03842_ net722 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a41o_1
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08881_ _04813_ _04814_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08194__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07832_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\]
+ net759 net1117 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07941__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11436__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ net1169 net874 team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\]
+ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__a21o_1
X_09502_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net1018 net539 _05443_
+ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08497__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07694_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\] net786
+ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09433_ _04648_ _04923_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14117__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11452__A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _05278_ _05281_ _05301_ _05193_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08315_ net1064 _04255_ _04256_ net1206 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09295_ net529 _03490_ _05144_ net607 vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10068__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1257_A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\]
+ net946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11598__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A1 _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ net845 _04103_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__o21a_4
XFILLER_0_15_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11556__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\] net733
+ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__a221o_1
XANTENNA__08421__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10007__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07059_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\]
+ net771 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__mux2_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_100_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
X_10070_ _02800_ _02811_ _05908_ _05913_ net1136 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__o41a_2
XANTENNA__11049__D net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10531__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13760_ clknet_leaf_133_wb_clk_i _01524_ _00125_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08488__A1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ _02931_ _05923_ _02829_ net688 vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12711_ net1398 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
X_13691_ clknet_leaf_27_wb_clk_i _01455_ _00056_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07160__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15042__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ net1355 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08147__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12036__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11244__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ net1381 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14312_ clknet_leaf_36_wb_clk_i _02076_ _00677_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\]
+ sky130_fd_sc_hd__dfrtp_1
X_11524_ _06409_ net617 net703 net696 vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08660__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14243_ clknet_leaf_25_wb_clk_i _02007_ _00608_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11455_ net495 net619 _06580_ net397 net1891 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11301__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] _06141_ vssd1 vssd1
+ vccd1 vccd1 _06231_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08948__C1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14174_ clknet_leaf_58_wb_clk_i _01938_ _00539_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[528\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08412__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ net507 net630 _06745_ net407 net2541 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a32o_1
X_13125_ net1274 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
X_10337_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] _06147_ _06149_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06974__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12921__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ net1407 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
X_10268_ _06107_ _06109_ _05979_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a21o_1
XANTENNA__13784__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1330 net1333 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__clkbuf_4
X_12007_ net1244 net657 net702 net473 vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__or4b_4
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1341 net1342 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__buf_4
Xfanout1352 net1359 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10199_ _04711_ _02774_ net672 vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__mux2_1
XANTENNA__10522__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1363 net1367 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__clkbuf_2
Xfanout1374 net1376 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__buf_4
Xfanout1385 net1386 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__buf_4
Xfanout1396 net1406 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08479__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ clknet_leaf_79_wb_clk_i _01722_ _00323_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12909_ net1291 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
XANTENNA__11483__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12368__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07151__A1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13889_ clknet_leaf_3_wb_clk_i _01653_ _00254_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12027__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10038__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08100__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08100_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[346\]
+ net765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\] net1119
+ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09080_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\]
+ net963 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\] net1067
+ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ net1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\]
+ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__or2_1
Xinput40 gpio_in[15] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput51 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput62 gpio_in[6] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11211__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\] vssd1
+ vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xinput73 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07197__A _03138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput84 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
Xhold813 team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\] vssd1
+ vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_1
XFILLER_0_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold824 team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\] vssd1
+ vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\] vssd1
+ vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07628__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold846 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\] vssd1
+ vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 team_03_WB.instance_to_wrap.core.register_file.registers_state\[429\] vssd1
+ vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ _05861_ net1948 net288 vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__mux2_1
Xhold868 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\] vssd1
+ vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\] vssd1
+ vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06965__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net1059 _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__nand2_1
XANTENNA__08520__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08167__B1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_A _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10989__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ net1200 _04805_ _04800_ net844 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12042__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15095__1476 vssd1 vssd1 vccd1 vccd1 _15095__1476/HI net1476 sky130_fd_sc_hd__conb_1
XANTENNA__10513__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1005_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ net1014 _02835_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1
+ vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__o21a_1
X_08795_ _04735_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__and2_1
XANTENNA__09116__C1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07746_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\] net726
+ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07660__A _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ net1106 _03615_ _03616_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout632_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1374_A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ net545 _04505_ _04478_ net561 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11182__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07693__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _04148_ _05287_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11332__D net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11777__A1 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_774 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09587__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09278_ _04893_ _05219_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ net1229 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\]
+ net955 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\] net916
+ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ net504 net625 _06687_ net413 net2172 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07602__C1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net632 _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nor2_1
XANTENNA__12741__A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06956__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ _03640_ _05961_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10912__D_N team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14930_ clknet_leaf_125_wb_clk_i _02685_ _01295_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10053_ net3 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1
+ vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ clknet_leaf_54_wb_clk_i _02625_ _01226_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07381__A1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11791__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ clknet_leaf_91_wb_clk_i _01576_ _00177_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\]
+ sky130_fd_sc_hd__dfrtp_1
X_14792_ clknet_leaf_32_wb_clk_i _02556_ _01157_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15199__1574 vssd1 vssd1 vccd1 vccd1 _15199__1574/HI net1574 sky130_fd_sc_hd__conb_1
XANTENNA__07570__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13743_ clknet_leaf_98_wb_clk_i _01507_ _00108_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_10955_ net510 net593 net264 net522 net1908 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07133__A1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12009__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10886_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[16\] net308 net685 vssd1
+ vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a21o_1
X_13674_ clknet_leaf_3_wb_clk_i _01438_ _00039_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07684__A2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11217__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12625_ net1312 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ net1303 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08605__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09830__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _06625_ net2566 net394 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__A3 net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ net1390 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XANTENNA__07841__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\] vssd1
+ vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14226_ clknet_leaf_105_wb_clk_i _01990_ _00591_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11438_ net280 net622 net704 net823 vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14157_ clknet_leaf_104_wb_clk_i _01921_ _00522_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\]
+ sky130_fd_sc_hd__dfrtp_1
X_11369_ net709 _06495_ net696 vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07295__S1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06947__B2 team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ net1323 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
X_14088_ clknet_leaf_27_wb_clk_i _01852_ _00453_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11267__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ net1388 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1160 team_03_WB.instance_to_wrap.core.decoder.inst\[21\] vssd1 vssd1 vccd1
+ vccd1 net1160 sky130_fd_sc_hd__clkbuf_8
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_2
Xfanout1182 net1197 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1193 net1196 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07600_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\]
+ net899 _03541_ net1149 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13482__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08580_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\] net919
+ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09649__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07531_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\] net795
+ net731 _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__o211a_1
XANTENNA__11456__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11206__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07462_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\]
+ net761 net1118 vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09201_ net605 _04071_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or2_1
XANTENNA__11208__A0 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07393_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[831\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[799\]
+ net768 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11759__A1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09132_ _04829_ net327 _05072_ _05073_ _04823_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08515__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07427__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ net1077 _05001_ _05004_ net844 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a31o_1
XANTENNA__10991__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08014_ net1107 _03954_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold610 team_03_WB.instance_to_wrap.core.register_file.registers_state\[567\] vssd1
+ vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\] vssd1
+ vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\] vssd1
+ vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\] vssd1
+ vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold654 team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\] vssd1
+ vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold665 net220 vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14305__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\] vssd1
+ vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold687 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\] vssd1
+ vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07060__B1 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 team_03_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net2282
+ sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _03756_ net661 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout582_A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\]
+ net958 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__mux2_1
X_09896_ net1120 _02804_ _05836_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__o211a_1
XANTENNA__09888__B1 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09870__A _05811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08847_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\]
+ net1008 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\] net1074
+ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__a221o_1
XANTENNA__07363__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout847_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08778_ net859 _04718_ _04719_ _04717_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a31o_1
X_07729_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\] net1143
+ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07115__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10740_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _05676_ net603 vssd1
+ vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__mux2_1
XANTENNA__11343__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__A1 net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10671_ _06311_ _05583_ _05563_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12410_ net1370 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ net1331 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
XANTENNA__08615__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12341_ net1263 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07823__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__B _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15060_ net1441 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12272_ net1417 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ clknet_leaf_28_wb_clk_i _01775_ _00376_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11786__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13567__A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06513_ net2653 net493 vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11154_ net1243 net828 _06478_ net669 vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__or4_1
X_10105_ team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] net672 vssd1 vssd1 vccd1
+ vccd1 _05949_ sky130_fd_sc_hd__nand2_1
X_11085_ _06620_ net2770 net424 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10036_ net21 net1034 _05907_ net1914 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__o22a_1
X_14913_ clknet_leaf_126_wb_clk_i _02668_ _01278_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11686__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08551__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14844_ clknet_leaf_55_wb_clk_i _02608_ _01209_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08396__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ clknet_leaf_60_wb_clk_i _02539_ _01140_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08303__B1 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ _06468_ net2351 net448 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13726_ clknet_leaf_78_wb_clk_i _01490_ _00091_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11253__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10938_ net296 net2432 net523 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10661__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ net685 _05833_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13657_ clknet_leaf_84_wb_clk_i _01421_ _00022_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11550__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ net1408 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08335__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15094__1475 vssd1 vssd1 vccd1 vccd1 _15094__1475/HI net1475 sky130_fd_sc_hd__conb_1
X_13588_ net1282 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10413__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08082__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ net1364 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14328__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13477__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ clknet_leaf_130_wb_clk_i _01973_ _00574_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15189_ net1570 vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07042__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout408 _06718_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14478__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout419 _06635_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
XANTENNA__07593__A1 net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06962_ net1157 _02901_ _02902_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__and3_1
X_09750_ _03727_ net588 vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__nor2_1
X_08701_ net1061 _04640_ _04641_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__or3_1
X_09681_ net582 _05501_ _05612_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__a31o_2
XANTENNA__11677__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06893_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] net1015 vssd1
+ vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08542__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\] net1204
+ vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11429__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08563_ net440 net432 _04503_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nor3_1
XANTENNA__09098__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07514_ _03451_ _03455_ _03454_ net1114 vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a2bb2o_1
X_08494_ net853 _04434_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07445_ net1106 _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08753__B net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A _06560_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\]
+ net894 net1122 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\] net1069
+ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11601__A0 _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1278_A team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1337_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09046_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\]
+ net988 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\] net942
+ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09022__A1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\] vssd1
+ vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07259__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold451 team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\] vssd1
+ vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_03_WB.instance_to_wrap.core.register_file.registers_state\[531\] vssd1
+ vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\] vssd1
+ vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07033__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold484 team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\] vssd1
+ vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold495 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\] vssd1
+ vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout964_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07584__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout920 net924 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11380__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 net932 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ _05878_ net1814 net292 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__mux2_1
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout953 net954 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_2
Xfanout964 net967 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_2
Xfanout975 net980 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout986 net987 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout997 net999 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
X_09879_ _05635_ _05813_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__o21ba_4
XANTENNA__11057__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\] vssd1
+ vssd1 vccd1 vccd1 net2724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\] vssd1
+ vssd1 vccd1 vccd1 net2735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\] vssd1
+ vssd1 vccd1 vccd1 net2746 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ _06611_ net2835 net373 vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__mux2_1
Xhold1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\] vssd1
+ vssd1 vccd1 vccd1 net2757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ net1370 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
Xhold1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\] vssd1
+ vssd1 vccd1 vccd1 net2768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[603\] vssd1
+ vssd1 vccd1 vccd1 net2779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10891__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09089__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _06679_ net482 net330 net2265 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14560_ clknet_leaf_1_wb_clk_i _02324_ _00925_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\]
+ sky130_fd_sc_hd__dfrtp_1
X_11772_ _06605_ net475 net338 net2669 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13511_ net1327 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
X_10723_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] net601 vssd1 vssd1 vccd1
+ vccd1 _06353_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14491_ clknet_leaf_30_wb_clk_i _02255_ _00856_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input93_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13442_ net1401 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10654_ net1246 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] net841 vssd1 vssd1 vccd1
+ vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ net1422 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ net1909 net535 net596 net590 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10946__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15112_ net1493 vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_2
XFILLER_0_134_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ net1306 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14620__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15043_ clknet_leaf_31_wb_clk_i _02763_ _01408_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12255_ net1374 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06911__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07024__B1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ net275 net2587 net493 vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__mux2_1
X_12186_ net1650 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ net2213 net420 _06644_ net519 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08119__A3 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ net832 _06414_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11123__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08838__B net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ net80 net79 net82 net81 vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14827_ clknet_leaf_31_wb_clk_i net1798 _01192_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ clknet_leaf_122_wb_clk_i _02522_ _01123_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08827__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13709_ clknet_leaf_105_wb_clk_i _01473_ _00074_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11831__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14689_ clknet_leaf_42_wb_clk_i _02453_ _01054_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07230_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07161_ _03075_ _03081_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\]
+ net876 _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09004__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__S0 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09555__A2 _05106_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07636__C net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07566__A1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11362__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ net540 _05741_ _05743_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07994_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\] net745
+ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o221a_1
XANTENNA__10570__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06945_ _02881_ _02886_ net818 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__mux2_1
X_09733_ _05673_ _05674_ _05668_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__a21o_1
XANTENNA__07318__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout378_A _06813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ _02814_ net1014 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__or2_2
X_09664_ _03170_ _04207_ net663 _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08615_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\] net921
+ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__a221o_1
X_09595_ net576 _05535_ _05536_ _04832_ _05534_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__a311o_1
XFILLER_0_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_71_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout545_A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08818__A1 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\] net996 net931
+ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07177__S0 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08477_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\] net928
+ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a221o_1
XANTENNA__11822__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__or3_1
XFILLER_0_17_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07359_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\] net1115
+ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _06200_ _06201_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] net677
+ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11050__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08703__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ net1239 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\]
+ net981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\] net928
+ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12040_ net1243 net653 _06463_ net468 vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__or4b_4
XFILLER_0_103_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold270 team_03_WB.instance_to_wrap.core.register_file.registers_state\[53\] vssd1
+ vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11889__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11349__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\] vssd1
+ vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\] vssd1
+ vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08754__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 net751 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__buf_4
Xfanout761 net766 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__buf_4
Xfanout772 net785 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07309__A1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13991_ clknet_leaf_64_wb_clk_i _01755_ _00356_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout783 net784 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_2
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11365__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15093__1474 vssd1 vssd1 vccd1 vccd1 _15093__1474/HI net1474 sky130_fd_sc_hd__conb_1
XFILLER_0_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12942_ net1336 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XANTENNA__11084__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ net1247 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13580__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07989__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14612_ clknet_leaf_91_wb_clk_i _02376_ _00977_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[966\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11824_ _06655_ net466 net328 net2241 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10616__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14543_ clknet_leaf_99_wb_clk_i _02307_ _00908_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11813__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ net646 _06580_ net458 net337 net2459 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a32o_1
XANTENNA__11304__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06906__B net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10706_ _06341_ _06342_ net604 vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ clknet_leaf_3_wb_clk_i _02238_ _00839_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11686_ _06728_ net387 net344 net1992 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ net1402 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10637_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] team_03_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ net840 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XANTENNA__08037__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10919__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10568_ net1797 net534 net595 _05878_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13356_ net1285 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
XANTENNA__09785__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12307_ net1264 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
X_10499_ net2229 net1028 net903 net1794 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
X_13287_ net1332 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15026_ clknet_leaf_33_wb_clk_i _02746_ _01391_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11259__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ net1639 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11344__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12169_ net1720 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08849__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A3 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11275__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07181__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ net1238 team_03_WB.instance_to_wrap.core.register_file.registers_state\[729\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\] net943
+ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__o221a_1
XANTENNA__13490__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _03566_ _05158_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08331_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[597\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14666__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09399__B _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11280__A1 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _04200_ _04201_ _04202_ _04203_ net855 net929 vssd1 vssd1 vccd1 vccd1 _04204_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07213_ net1106 _03153_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08193_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\]
+ net947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\] net913
+ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07144_ net733 _03082_ _03083_ _03084_ _03085_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a32o_1
XANTENNA__07787__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07331__S0 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08984__B1 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12045__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\]
+ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__B1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1035_A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07539__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09862__B _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10543__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11886__A3 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _03916_ _03918_ net1159 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__o21a_1
X_09716_ _04832_ _05548_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__or2_1
X_06928_ net1147 net1114 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_4
XFILLER_0_138_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09700__A2 _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ net1109 _02804_ net539 _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06859_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] vssd1 vssd1 vccd1
+ vccd1 _02801_ sky130_fd_sc_hd__and3b_2
XANTENNA__07711__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout927_A net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07172__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08494__A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ net573 _05399_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__nand2_1
X_08529_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\]
+ net970 net1071 vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11540_ net502 net623 _06650_ net487 net1869 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__a32o_1
XANTENNA__07475__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11351__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ net656 _06596_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09216__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11023__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ _06064_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__xnor2_1
X_13210_ net1365 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
X_14190_ clknet_leaf_70_wb_clk_i _01954_ _00555_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07778__A1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ _06104_ _06089_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__nand2b_1
X_13141_ net1262 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10782__B1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ net1427 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
X_10284_ _06125_ _06123_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nand2b_1
XANTENNA_input56_A gpio_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12023_ net634 _06585_ net472 net368 net2195 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__a32o_1
XANTENNA__08727__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10534__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14539__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11095__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _02993_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_4
X_13974_ clknet_leaf_86_wb_clk_i _01738_ _00339_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[328\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12925_ net1381 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XANTENNA__07702__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12039__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ net1368 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11807_ net2478 _06632_ net333 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12787_ net1265 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14526_ clknet_leaf_58_wb_clk_i _02290_ _00891_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[880\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07466__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11262__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11261__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ net593 net264 net475 _06808_ net1887 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a32o_1
XANTENNA__10158__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14457_ clknet_leaf_111_wb_clk_i _02221_ _00822_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09207__A1 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ net2034 net265 net349 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11014__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ net1424 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XANTENNA__07748__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__A2 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14069__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14388_ clknet_leaf_91_wb_clk_i _02152_ _00753_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11565__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13339_ net1286 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XANTENNA__10174__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09963__A _03723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08981__A3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\] net781
+ _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__a21o_1
X_15009_ clknet_leaf_23_wb_clk_i net57 _01374_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08880_ net560 _04770_ net540 _04819_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10902__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[13\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08194__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ _03769_ _03770_ _03772_ net1115 vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__o22a_1
XANTENNA__07941__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11209__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11436__C net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__or3_1
X_09501_ _03823_ _04444_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07693_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\] net758
+ net1011 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12829__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09432_ _05372_ _05373_ net556 vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10994__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _05291_ _05303_ _05304_ _05288_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\]
+ net983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\] net1217
+ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09294_ _05226_ _05228_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08245_ net855 _04183_ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09857__B _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout410_A _06717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1152_A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout508_A net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ net1199 _04110_ _04117_ net845 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__o211ai_1
X_15092__1473 vssd1 vssd1 vccd1 vccd1 _15092__1473/HI net1473 sky130_fd_sc_hd__conb_1
XANTENNA__09749__A2 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11556__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\] net778 net733
+ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__a221o_1
XANTENNA__08957__B1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07058_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\]
+ net771 vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__mux2_1
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_98_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__11908__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XANTENNA__10516__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A2 _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10819__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _06550_ net2313 net522 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__B2 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ net1419 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13690_ clknet_leaf_20_wb_clk_i _01454_ _00055_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12641_ net1288 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11244__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ net1347 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XANTENNA__08645__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07999__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ clknet_leaf_65_wb_clk_i _02075_ _00676_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11789__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11523_ net2106 net488 _06780_ net506 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14242_ clknet_leaf_131_wb_clk_i _02006_ _00607_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\]
+ sky130_fd_sc_hd__dfrtp_1
X_11454_ net502 net621 _06579_ net398 net1946 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10204__C1 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net285 _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__and2_1
X_14173_ clknet_leaf_68_wb_clk_i _01937_ _00538_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\]
+ sky130_fd_sc_hd__dfrtp_1
X_11385_ net716 net269 net699 vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06959__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13124_ net1307 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
X_10336_ _06172_ _06173_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] net675
+ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__o2bb2a_1
X_15188__1569 vssd1 vssd1 vccd1 vccd1 _15188__1569/HI net1569 sky130_fd_sc_hd__conb_1
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10267_ _05979_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13055_ net1375 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XANTENNA__08176__A1 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1320 net1335 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__buf_4
X_12006_ _06557_ net2584 net451 vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__mux2_1
Xfanout1331 net1332 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__buf_4
X_10198_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] net659 _06038_ _02889_
+ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__o211a_1
Xfanout1342 net1359 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__buf_2
XANTENNA__07384__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1353 net1358 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__buf_4
Xfanout1364 net1367 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__buf_4
XFILLER_0_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1375 net1376 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1386 net1387 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__clkbuf_4
Xfanout1397 net1406 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__buf_4
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13957_ clknet_leaf_109_wb_clk_i _01721_ _00322_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ net1303 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
XANTENNA__07687__B1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ clknet_leaf_133_wb_clk_i _01652_ _00253_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_128_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12839_ net1399 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10169__A _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10038__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08862__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08100__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__C_N net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14509_ clknet_leaf_106_wb_clk_i _02273_ _00874_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08030_ net811 _03967_ _03968_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__o22ai_2
XANTENNA__14704__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 gpio_in[16] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput52 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput63 gpio_in[7] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
Xhold803 team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\] vssd1
+ vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
Xhold814 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\] vssd1
+ vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput85 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
Xhold825 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\] vssd1
+ vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xinput96 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold836 team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\] vssd1
+ vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\] vssd1
+ vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold858 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\] vssd1
+ vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09039__S0 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ _05852_ _05858_ _05082_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__or3b_1
Xhold869 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\] vssd1
+ vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_08932_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\]
+ net972 net1070 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08167__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10989__D net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08863_ net1063 _04801_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a21o_1
XANTENNA__07914__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__S1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07814_ net718 _03739_ _03748_ _03755_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__06865__C_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08794_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[706\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\] net921
+ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__a221o_1
XANTENNA__09116__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ net726 _03683_ _03684_ _03685_ _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07127__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout458_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07678__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ net1152 _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__or2_1
XANTENNA__11474__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09415_ _04416_ _04533_ net551 vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__mux2_1
XANTENNA__08475__C _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12018__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1367_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09346_ _04148_ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08627__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _03759_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11402__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14384__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08228_ _04166_ _04169_ net1077 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09052__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08159_ net1055 _04098_ _04099_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__or3_1
XANTENNA__10737__B1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11170_ net716 _06503_ net694 vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__or3_1
XFILLER_0_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ _05962_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10542__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ net4 net1033 net907 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1
+ vccd1 vccd1 _02679_ sky130_fd_sc_hd__o22a_1
XANTENNA__11357__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11701__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ clknet_leaf_41_wb_clk_i net1990 _01225_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ clknet_leaf_113_wb_clk_i _01575_ _00176_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791_ clknet_leaf_31_wb_clk_i _02555_ _01156_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11373__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ clknet_leaf_69_wb_clk_i _01506_ _00107_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11465__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ net829 _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13673_ clknet_leaf_77_wb_clk_i _01437_ _00038_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10885_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[16\] net306 vssd1
+ vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ net1427 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
XANTENNA__14727__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__S1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08618__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11768__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08094__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12555_ net1257 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11312__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11506_ _06624_ net2840 net394 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__mux2_1
XANTENNA__10440__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07841__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12486_ net1412 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ clknet_leaf_96_wb_clk_i _01989_ _00590_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09189__A3 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ net2797 net400 _06758_ net506 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08397__A1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ clknet_leaf_5_wb_clk_i _01920_ _00521_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06930__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11368_ net499 net619 _06736_ net405 net1894 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06947__A2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ net1264 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
X_10319_ net282 _06159_ net675 vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10452__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ clknet_leaf_68_wb_clk_i _01851_ _00452_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08149__A1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ net1038 _06449_ net649 _06463_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__or4_4
XANTENNA__11267__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ net1283 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09897__A1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1150 team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1 vccd1
+ vccd1 net1150 sky130_fd_sc_hd__buf_4
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11982__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1161 net1163 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1172 net1178 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_2
Xfanout1183 net1197 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10900__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1194 net1195 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__buf_2
XANTENNA__07761__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09649__A1 _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15091__1472 vssd1 vssd1 vccd1 vccd1 _15091__1472/HI net1472 sky130_fd_sc_hd__conb_1
X_14989_ clknet_leaf_41_wb_clk_i net37 _01354_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__07109__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11283__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07755__S0 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07461_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\] net1143
+ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ _02954_ _05107_ _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07392_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09131_ net584 _02953_ net581 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__and3_2
XFILLER_0_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08085__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11222__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09062_ net926 _05003_ _05002_ net1215 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08013_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\]
+ net760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\] net728
+ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09034__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold600 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\] vssd1
+ vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\] vssd1
+ vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08388__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\] vssd1
+ vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10065__C net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold633 team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\] vssd1
+ vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold644 team_03_WB.instance_to_wrap.core.register_file.registers_state\[755\] vssd1
+ vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold655 net190 vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\] vssd1
+ vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold677 team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\] vssd1
+ vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 net160 vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11458__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09964_ _05886_ net1913 net292 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12053__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold699 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\] vssd1
+ vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15032__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1115_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08915_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\]
+ net958 vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__mux2_1
XANTENNA__07374__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _04031_ _04323_ net539 vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__or3_1
XANTENNA__09888__A1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10498__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__B1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08846_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\]
+ net1008 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\] net1207
+ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a221o_1
XANTENNA__08560__A1 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout742_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\] net921
+ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ net1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\] net1120
+ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__o221a_1
XANTENNA__11447__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08312__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11998__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07659_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] net1012 _03107_ vssd1
+ vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__a21o_2
XANTENNA__11343__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187__1568 vssd1 vssd1 vccd1 vccd1 _15187__1568/HI net1568 sky130_fd_sc_hd__conb_1
XANTENNA__07520__C1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ _05583_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09902__D_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ _05246_ _05250_ _05269_ _05244_ _05241_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__a311o_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12340_ net1304 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07823__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10971__S net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ net1407 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__inv_2
XANTENNA__12752__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14010_ clknet_leaf_21_wb_clk_i _01774_ _00375_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\]
+ sky130_fd_sc_hd__dfrtp_1
X_11222_ net270 net2578 net490 vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XANTENNA__09671__S0 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11153_ net494 net646 _06653_ net417 net2091 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ _02811_ _02816_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a211o_1
X_11084_ net827 net274 vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__and2_1
XANTENNA__11135__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ clknet_leaf_38_wb_clk_i _00006_ _01277_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10035_ net22 net1033 net907 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1
+ vccd1 vccd1 _02696_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ clknet_leaf_54_wb_clk_i net1933 _01208_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output125_A net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06909__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14774_ clknet_leaf_56_wb_clk_i _02538_ _01139_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__C net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ _06453_ net2716 net448 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13725_ clknet_leaf_66_wb_clk_i _01489_ _00090_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10937_ net686 _06521_ _06522_ _06520_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__o31a_4
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ clknet_leaf_11_wb_clk_i _01420_ _00021_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06925__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10868_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[19\] net308 net685 vssd1
+ vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09301__A _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ net1377 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09803__A1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ net1280 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10949__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[30\] net307 _06407_ net692
+ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12538_ net1365 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11977__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09955__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12469_ net1261 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09567__B1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ clknet_leaf_132_wb_clk_i _01972_ _00573_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08351__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1569 vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_2
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11374__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07042__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ clknet_leaf_28_wb_clk_i _01903_ _00504_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[493\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10182__A team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout409 net410 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09971__A _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06961_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[389\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[261\]
+ net770 net1121 vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__mux4_1
XANTENNA__13493__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\]
+ net977 net1073 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux4_1
X_09680_ _05621_ _05616_ _05620_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__or3b_1
XFILLER_0_20_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06892_ _02816_ _02830_ _02833_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nor3_1
XFILLER_0_20_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08631_ net859 _04571_ _04572_ _04570_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08562_ _04503_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07513_ net1124 _03453_ net1160 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08493_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\]
+ net988 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\] net942
+ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o221a_1
X_07444_ net1151 _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09211__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10357__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ net1090 net893 team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\]
+ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1065_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\]
+ net949 net1069 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09045_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\] net1006
+ net926 _04986_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__o211a_1
XANTENNA__10955__A3 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07281__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1232_A net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold430 team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\] vssd1
+ vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\] vssd1
+ vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 team_03_WB.instance_to_wrap.CPU_DAT_I\[7\] vssd1 vssd1 vccd1 vccd1 net2036
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14422__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold463 team_03_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1 net2047
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11188__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 net108 vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10092__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08230__B1 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\] vssd1
+ vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 team_03_WB.instance_to_wrap.ADR_I\[1\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout910 net912 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout921 net924 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09947_ _03389_ net660 vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__nor2_1
Xfanout932 net936 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_4
Xfanout943 net944 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
Xfanout954 net968 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout957_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 net980 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14572__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ net358 _05404_ _05815_ _05817_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a2111o_1
Xfanout987 net992 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_2
Xhold1130 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\] vssd1
+ vssd1 vccd1 vccd1 net2714 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
Xhold1141 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\] vssd1
+ vssd1 vccd1 vccd1 net2725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\] vssd1
+ vssd1 vccd1 vccd1 net2736 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ _04080_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__nor2_1
Xhold1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\] vssd1
+ vssd1 vccd1 vccd1 net2747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\] vssd1
+ vssd1 vccd1 vccd1 net2758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\] vssd1
+ vssd1 vccd1 vccd1 net2769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\] vssd1
+ vssd1 vccd1 vccd1 net2780 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ _06678_ net477 net329 net2029 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10891__A2 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__S1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11771_ net654 _06604_ net475 net338 net2103 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a32o_1
XANTENNA__07639__A3 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ net1327 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10722_ net1731 net531 net528 _06352_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08436__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09685__A1_N net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490_ clknet_leaf_22_wb_clk_i _02254_ _00855_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[844\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ net1401 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ net1245 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] net841 vssd1 vssd1 vccd1
+ vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13372_ net1423 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XANTENNA_input86_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ net1871 net536 net597 _02888_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11797__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15111_ net1492 vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_2
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ net1297 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15090__1471 vssd1 vssd1 vccd1 vccd1 _15090__1471/HI net1471 sky130_fd_sc_hd__conb_1
XFILLER_0_106_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09549__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15042_ clknet_leaf_32_wb_clk_i _02762_ _01407_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dfrtp_1
X_12254_ net1384 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09644__S0 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11205_ net277 net2412 net493 vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07024__A1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ net1629 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11136_ net276 net657 net707 net698 vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11659__A1 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _06611_ net2781 net421 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XANTENNA__08524__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ _05892_ _05893_ _05894_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07742__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14826_ clknet_leaf_32_wb_clk_i net2006 _01191_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09730__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14757_ clknet_leaf_123_wb_clk_i _02521_ _01122_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12657__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ net636 _06746_ net475 net371 net2141 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11561__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ clknet_leaf_9_wb_clk_i _01472_ _00073_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11831__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14688_ clknet_leaf_42_wb_clk_i _02452_ _01053_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13639_ net1424 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XANTENNA__10177__A _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07160_ net814 _03091_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11595__A0 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14445__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13488__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\]
+ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11500__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08438__S1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08212__B1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15186__1567 vssd1 vssd1 vccd1 vccd1 _15186__1567/HI net1567 sky130_fd_sc_hd__conb_1
X_09801_ _03490_ _04592_ net665 _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07993_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\] net735
+ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _02953_ net577 _05442_ net360 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a31o_1
X_06944_ _02882_ _02883_ _02885_ _02884_ net747 net809 vssd1 vssd1 vccd1 vccd1 _02886_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09663_ net541 _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06875_ _02794_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] _02805_
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a2111oi_2
XANTENNA_fanout273_A _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08614_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\] net938
+ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ net570 _05407_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout440_A _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07177__S1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11822__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11190__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07427_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\] net787
+ net1011 _03368_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout705_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07358_ net1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[668\] net786 net737
+ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__o221a_1
XANTENNA__11586__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08451__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11050__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\]
+ net778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\] net748
+ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11410__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13812__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ _04964_ _04969_ net870 vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__mux2_1
XANTENNA__14938__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07827__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11338__B1 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold260 net226 vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11889__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold271 team_03_WB.instance_to_wrap.core.register_file.registers_state\[564\] vssd1
+ vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11349__C net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10010__A0 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold282 team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\] vssd1
+ vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold293 team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\] vssd1
+ vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
Xfanout751 _02852_ vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
Xfanout762 net765 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
X_13990_ clknet_leaf_78_wb_clk_i _01754_ _00355_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout773 net776 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
Xfanout784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__clkbuf_4
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_2
XANTENNA__11365__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ net1291 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XANTENNA__10313__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12872_ net1285 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
X_14611_ clknet_leaf_115_wb_clk_i _02375_ _00976_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_90_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11823_ net646 _06653_ net457 net328 net1911 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11381__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ clknet_leaf_76_wb_clk_i _02306_ _00907_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11754_ net651 _06579_ net461 net340 net1985 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a32o_1
XANTENNA__11813__A1 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__A2 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10705_ team_03_WB.instance_to_wrap.core.pc.current_pc\[26\] _06315_ vssd1 vssd1
+ vccd1 vccd1 _06342_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ clknet_leaf_58_wb_clk_i _02237_ _00838_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11685_ _06727_ net388 net347 net2165 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13424_ net1400 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10636_ team_03_WB.instance_to_wrap.core.decoder.inst\[25\] team_03_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ net842 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XANTENNA__11577__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_107_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07245__A1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ net1286 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
X_10567_ net1858 net534 net595 _05877_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__A3 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06922__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ net1410 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286_ net1332 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XANTENNA__11329__A0 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498_ net133 net1027 net903 net2070 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15025_ clknet_leaf_31_wb_clk_i _02745_ _01390_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12237_ net1745 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11259__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10001__A0 _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08745__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ net1743 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10552__A1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07953__C1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11119_ _06633_ net2774 net423 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__mux2_1
XANTENNA__06885__A_N _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12099_ _06796_ net479 net446 net2115 vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09026__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11501__A0 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11990__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07181__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ clknet_leaf_56_wb_clk_i net1704 _01174_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11291__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08330_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11804__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07484__A1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08261_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1010\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11280__A2 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07212_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\] net724
+ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08192_ _04128_ _04133_ net867 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07143_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\]
+ net879 net1149 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__o211a_1
XANTENNA__11230__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__S1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08984__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\]
+ net798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[354\] net1146
+ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_105_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10791__A1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__A1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout390_A net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout488_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12061__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\]
+ net900 _03917_ net1147 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__o311a_1
XFILLER_0_138_1414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09715_ _04777_ _05650_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a21oi_2
X_06927_ net1116 net1151 vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nor2_8
XFILLER_0_39_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout655_A _06457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1397_A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09646_ _03428_ _04295_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06858_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__nand4b_4
XANTENNA__07172__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09577_ _05315_ _05431_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11405__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08528_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\]
+ net972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o221a_1
XANTENNA__09464__A2 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__A3 _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07475__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08459_ net845 _04400_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14760__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11470_ net496 net620 _06595_ net397 net2471 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10421_ _06012_ _06014_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__nand2_1
XANTENNA__07227__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11023__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ net1323 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10352_ team_03_WB.instance_to_wrap.core.pc.current_pc\[23\] _06147_ vssd1 vssd1
+ vccd1 vccd1 _06186_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ net1388 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
X_10283_ _05973_ _06124_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__nand2_1
XANTENNA__08727__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09545__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _06766_ net466 net366 net2335 vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__a22o_1
XANTENNA_input49_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11731__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14140__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _03024_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_4
Xfanout581 _02992_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
Xfanout592 _02951_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__buf_4
XANTENNA__11095__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ clknet_leaf_88_wb_clk_i _01737_ _00338_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09152__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ net1342 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07702__A2 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14290__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12855_ net1418 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11315__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ net2491 net263 net333 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12786_ net1420 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14525_ clknet_leaf_66_wb_clk_i _02289_ _00890_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07466__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15185__1566 vssd1 vssd1 vccd1 vccd1 _15185__1566/HI net1566 sky130_fd_sc_hd__conb_1
XANTENNA__11262__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ net1939 net269 net342 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07561__S1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14456_ clknet_leaf_10_wb_clk_i _02220_ _00821_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11668_ net1999 _06629_ net349 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
X_13407_ net1326 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XANTENNA__07218__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11014__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ net1604 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] net837 vssd1 vssd1 vccd1
+ vccd1 _02509_ sky130_fd_sc_hd__mux2_1
X_14387_ clknet_leaf_110_wb_clk_i _02151_ _00752_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\]
+ sky130_fd_sc_hd__dfrtp_1
X_11599_ _06518_ net2460 net454 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07769__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ net1292 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10174__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11985__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11970__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ net1263 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XANTENNA__12670__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15008_ clknet_leaf_124_wb_clk_i net56 _01373_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07764__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07077__S0 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11722__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ net1166 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\]
+ net872 _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\]
+ net888 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__or3_1
XANTENNA__14633__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11436__D net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07692_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\] net786
+ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07154__B1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _05013_ _05070_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13006__A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09362_ _05283_ _05289_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__nand2_1
XANTENNA__14783__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\]
+ net983 vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08654__B1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _05222_ _05233_ _05234_ _05220_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_35_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15221__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08244_ net850 _04184_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06843__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07209__A1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _04114_ _04116_ net1077 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout403_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1145_A team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08957__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07126_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\] net778
+ net749 _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10084__B _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11961__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07057_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\]
+ net772 net1122 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__mux4_1
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1312_A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14163__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__11908__B net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ net1139 net1017 net682 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10819__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ _06547_ _06548_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__a21oi_4
XANTENNA__08342__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _03314_ _04415_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or2_1
XANTENNA__10091__A_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12640_ net1379 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07448__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ net1364 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XANTENNA__08645__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ clknet_leaf_79_wb_clk_i _02074_ _00675_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07849__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _06405_ net631 net705 net699 vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14241_ clknet_leaf_0_wb_clk_i _02005_ _00606_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ net2806 net397 _06765_ net501 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08948__A1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14506__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _06070_ _06079_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__xnor2_1
X_14172_ clknet_leaf_128_wb_clk_i _01936_ _00537_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[526\]
+ sky130_fd_sc_hd__dfrtp_1
X_11384_ net513 net638 _06744_ net407 net2186 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a32o_1
XANTENNA__10755__A1 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13123_ net1262 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
X_10335_ net282 _06151_ _06169_ net675 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__o31a_1
XANTENNA__07620__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13054_ net1378 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
X_10266_ _03528_ _05978_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11704__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1310 net1317 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ net267 net2462 net451 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__mux2_1
Xfanout1321 net1335 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1332 net1333 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__buf_4
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10197_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] net659 _06038_ vssd1
+ vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__o21ai_1
Xfanout1343 net1345 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__buf_4
XANTENNA__07384__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1354 net1358 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__buf_2
Xfanout1365 net1367 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__buf_4
Xfanout1376 net1380 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__clkbuf_4
Xfanout1387 net1433 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__clkbuf_4
Xfanout1398 net1399 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__buf_4
XANTENNA__09125__A1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07136__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ clknet_leaf_15_wb_clk_i _01720_ _00321_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06928__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09676__A2 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07523__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ net1271 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_13887_ clknet_leaf_122_wb_clk_i _01651_ _00252_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11483__A2 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07151__A3 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ net1416 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10169__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12769_ net1276 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14508_ clknet_leaf_5_wb_clk_i _02272_ _00873_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
XFILLER_0_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14439_ clknet_leaf_63_wb_clk_i _02203_ _00804_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14186__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput42 gpio_in[17] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput64 gpio_in[8] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
Xinput75 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_1
Xhold804 team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\] vssd1
+ vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
Xhold815 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\] vssd1
+ vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\] vssd1
+ vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
Xhold837 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11943__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold848 team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\] vssd1
+ vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09980_ _03103_ net2061 net294 vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__mux2_1
Xhold859 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\] vssd1
+ vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09039__S1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08931_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09364__A1 _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ net1216 _04802_ _04803_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08572__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ net820 _03754_ net723 vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\] net938
+ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__a221o_1
XANTENNA__09116__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07744_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\]
+ net888 net1118 vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_36_1503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09214__A _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\]
+ net759 net1115 vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__mux4_1
XANTENNA__11474__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ net325 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1095_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _03137_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08627__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout520_A _06448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1262_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10434__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07669__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _03244_ _03790_ _05145_ net607 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ net1059 _04167_ _04168_ net1206 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__a211o_1
XANTENNA__07388__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09052__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\]
+ net950 net1066 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10198__C1 _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11934__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07109_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\] net731
+ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__a221oi_1
XANTENNA__07602__A1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08089_ _04029_ _04030_ net608 vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__mux2_2
XANTENNA__10823__A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09095__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _03640_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08789__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ net5 net1032 net906 net2862 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__o22a_1
XANTENNA__11357__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15184__1565 vssd1 vssd1 vccd1 vccd1 _15184__1565/HI net1565 sky130_fd_sc_hd__conb_1
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09107__A1 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ clknet_leaf_101_wb_clk_i _01574_ _00175_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ clknet_leaf_32_wb_clk_i _02554_ _01155_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08315__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ clknet_leaf_104_wb_clk_i _01505_ _00106_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11465__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07570__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _06533_ _06534_ _06535_ _06399_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__o211a_2
XFILLER_0_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ clknet_leaf_18_wb_clk_i _01436_ _00037_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10884_ net508 net593 _06479_ net522 net1769 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12623_ net1389 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08618__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12485__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12554_ net1258 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10976__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09830__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06623_ net2691 net395 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__mux2_1
XANTENNA__06914__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12485_ net1276 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14224_ clknet_leaf_81_wb_clk_i _01988_ _00589_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[578\]
+ sky130_fd_sc_hd__dfrtp_1
X_11436_ _06405_ net631 net705 net826 vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10728__A1 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14155_ clknet_leaf_17_wb_clk_i _01919_ _00520_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07054__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ net710 _06491_ net695 vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__and3_1
XANTENNA__06930__B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ net1420 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
X_10318_ _06153_ _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14086_ clknet_leaf_79_wb_clk_i _01850_ _00451_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\]
+ sky130_fd_sc_hd__dfrtp_1
X_11298_ net517 net642 _06716_ net416 net2336 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a32o_1
XANTENNA__10452__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ net1318 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
X_10249_ _03426_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11267__C net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11153__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__clkbuf_8
Xfanout1151 net1152 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1162 net1163 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_2
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1173 net1174 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10900__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1184 net1185 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_2
Xfanout1195 net1196 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07109__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14988_ clknet_leaf_107_wb_clk_i net36 _01353_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12102__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11283__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11456__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ clknet_leaf_113_wb_clk_i _01703_ _00304_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09969__A _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\] net1118
+ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o221a_1
XANTENNA__07755__S1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07391_ net818 _03324_ _03327_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__o22ai_1
XANTENNA__11503__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09130_ _04895_ _04956_ _05014_ _05071_ net559 net568 vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11759__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__A1 net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09282__B1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__A3 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09061_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\]
+ net986 vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08012_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\]
+ net760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\] net742
+ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold601 team_03_WB.instance_to_wrap.core.register_file.registers_state\[313\] vssd1
+ vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold612 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\] vssd1
+ vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold623 team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\] vssd1
+ vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07045__C1 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10065__D team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\] vssd1
+ vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 net132 vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold656 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\] vssd1
+ vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07596__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\] vssd1
+ vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08793__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _03723_ net660 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\] vssd1
+ vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 _02602_ vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08914_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\]
+ net958 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__mux2_1
X_09894_ _04031_ _04323_ net663 _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1010_A _04085_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09888__A2 _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _04783_ _04786_ net864 vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11695__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__S0 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15059__1440 vssd1 vssd1 vccd1 vccd1 _15059__1440/HI net1440 sky130_fd_sc_hd__conb_1
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08776_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\] net938
+ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__a221o_1
X_07727_ _03663_ _03668_ net1133 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10655__A0 team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07658_ _03585_ _03586_ _03599_ net720 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__a22o_4
XFILLER_0_95_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08783__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07520__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout902_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07589_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\] net782
+ net749 _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ _05246_ _05250_ _05269_ _05244_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ _05012_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12270_ net1338 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08722__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11907__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ net2365 net492 _06682_ net507 vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XANTENNA__07587__A0 _03526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07338__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ net703 net273 net695 vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__and3_1
XANTENNA__07051__A2 _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ net680 net284 vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
X_11083_ _06619_ net2310 net421 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__mux2_1
XANTENNA__11135__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ clknet_leaf_39_wb_clk_i _00005_ _01276_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10034_ net23 net1034 _05907_ net2860 vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__o22a_1
XANTENNA__11686__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10894__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ clknet_leaf_55_wb_clk_i _02606_ _01207_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08169__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14773_ clknet_leaf_55_wb_clk_i _02537_ _01138_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11985_ net274 net2497 net449 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__mux2_1
XANTENNA__08839__B1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__D net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__A0 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13724_ clknet_leaf_118_wb_clk_i _01488_ _00089_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\] net313 net311 net321
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__and4_1
XFILLER_0_131_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10867_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[19\] net306 vssd1
+ vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__and2_1
X_13655_ clknet_leaf_72_wb_clk_i _01419_ _00020_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11323__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ net1385 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
X_13586_ net1336 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ net313 net311 net322 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09803__A2 _05403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12537_ net1354 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12943__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12468_ net1304 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11419_ net298 net2559 net402 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__mux2_1
X_14207_ clknet_leaf_117_wb_clk_i _01971_ _00572_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11559__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15187_ net1568 vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_2
X_12399_ net1407 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11374__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14138_ clknet_leaf_23_wb_clk_i _01902_ _00503_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10182__B _02819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09971__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\] net1121
+ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__a221o_1
X_14069_ clknet_leaf_87_wb_clk_i _01833_ _00434_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11677__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ _02799_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__nand2_1
X_08630_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\] net922
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07750__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ net845 _04502_ _04491_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10637__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07512_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\]
+ net775 net1124 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08492_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\]
+ net988 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\] net926
+ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__o221a_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07443_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\]
+ net756 net1116 vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11233__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\]
+ net878 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183__1564 vssd1 vssd1 vccd1 vccd1 _15183__1564/HI net1564 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09113_ _05049_ _05054_ net871 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__mux2_1
XANTENNA__07012__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1058_A _02790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09044_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\] net988
+ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__or2_1
XANTENNA__07947__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09007__B1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06851__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold420 team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\] vssd1
+ vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold431 net186 vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1225_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\] vssd1
+ vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 team_03_WB.instance_to_wrap.CPU_DAT_I\[30\] vssd1 vssd1 vccd1 vccd1 net2037
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08766__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold464 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\] vssd1
+ vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11188__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07033__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold475 _02617_ vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold486 team_03_WB.instance_to_wrap.ADR_I\[8\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout685_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 _02604_ vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__buf_2
XANTENNA__09881__B _05811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09946_ _05877_ net2239 net292 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 net936 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_4
XANTENNA__14717__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net957 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_4
XANTENNA__07682__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__clkbuf_4
Xfanout977 net979 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__clkbuf_4
Xhold1120 team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\] vssd1
+ vssd1 vccd1 vccd1 net2704 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout852_A _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _03604_ _05069_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__o21a_1
Xfanout988 net992 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\] vssd1
+ vssd1 vccd1 vccd1 net2715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 net1010 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_4
XANTENNA__11408__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1142 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\] vssd1
+ vssd1 vccd1 vccd1 net2726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__B1 _06472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _04769_ _04768_ _04754_ _04748_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a2bb2o_4
Xhold1153 team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\] vssd1
+ vssd1 vccd1 vccd1 net2737 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\] vssd1
+ vssd1 vccd1 vccd1 net2748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\] vssd1
+ vssd1 vccd1 vccd1 net2759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\] vssd1
+ vssd1 vccd1 vccd1 net2770 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13741__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08759_ net1060 _04697_ _04700_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__a21oi_1
Xhold1197 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\] vssd1
+ vssd1 vccd1 vccd1 net2781 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10891__A3 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11770_ net653 _06603_ net469 net339 net2237 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12093__A2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10721_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] _05623_ net601 vssd1
+ vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13440_ net1401 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
X_10652_ net1241 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\] net839 vssd1 vssd1 vccd1
+ vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XANTENNA__09246__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ net1324 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ net1676 net538 net599 _02921_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12322_ net1374 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
X_15110_ net1491 vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_2
XFILLER_0_84_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10800__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input79_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15041_ clknet_leaf_31_wb_clk_i _02761_ _01406_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11379__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ net1382 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11356__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09013__A3 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ net278 net2514 net490 vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__mux2_1
XANTENNA__08757__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__S0 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ net1628 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ net503 net651 _06643_ net417 net1875 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08509__C1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ net827 net280 vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11318__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__C_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ net71 net70 net73 net72 vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ clknet_leaf_41_wb_clk_i net1784 _01190_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12938__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ clknet_leaf_15_wb_clk_i _02520_ _01121_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11968_ net633 _06745_ net474 net372 net2344 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09312__A _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ clknet_leaf_46_wb_clk_i _01471_ _00072_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11292__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07496__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[10\] net309 net688 vssd1
+ vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a21oi_1
X_14687_ clknet_leaf_42_wb_clk_i _02451_ _01052_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ net636 _06708_ net476 net380 net2145 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13638_ net1424 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10177__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09788__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13569_ net1313 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07799__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08996__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07090_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\]
+ net876 _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11289__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ net542 _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__nand2_1
X_07992_ net1132 _03933_ net722 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10570__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07971__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06943_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\]
+ net773 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__mux2_1
X_09731_ net585 _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11228__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ _03170_ _04207_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__or2_1
X_06874_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ _02794_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__or3_1
XANTENNA__07723__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ _04553_ _04554_ net854 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o21a_1
XANTENNA__07007__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ net566 _05415_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__nand2_1
XANTENNA__12848__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_A _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08544_ net1056 _04484_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__or3_1
XANTENNA__06846__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__A2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09222__A _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ net437 net429 _04415_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or3_2
XFILLER_0_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12059__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1175_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\]
+ net886 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11190__C net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07239__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\]
+ net759 vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout600_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1342_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07677__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08987__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ net1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\]
+ net778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\] net733
+ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09027_ net1213 _04967_ _04968_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11338__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold250 team_03_WB.instance_to_wrap.core.register_file.registers_state\[404\] vssd1
+ vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold261 net126 vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\] vssd1
+ vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11349__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold283 team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\] vssd1
+ vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 net222 vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08754__A2 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net735 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09929_ _03277_ net660 vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nor2_1
Xfanout752 net755 vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10550__B net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout763 net765 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout774 net776 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_4
Xfanout785 _02851_ vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_6
XANTENNA__09703__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout796 net799 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_2
X_12940_ net1303 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
XANTENNA__08062__S0 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11365__C net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__C1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12871_ net1398 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ clknet_leaf_100_wb_clk_i _02374_ _00975_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\]
+ sky130_fd_sc_hd__dfstp_1
X_11822_ net646 _06652_ net456 net328 net2083 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08447__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__A1 _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__B net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11753_ _06578_ net463 net337 net2384 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
XANTENNA__11274__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ clknet_leaf_106_wb_clk_i _02305_ _00906_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ _05933_ _06310_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__nor2_1
XANTENNA__10709__C net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ clknet_leaf_34_wb_clk_i _02236_ _00837_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _06726_ net390 net346 net2227 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ net1403 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
X_10635_ team_03_WB.instance_to_wrap.core.decoder.inst\[26\] team_03_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ net842 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11601__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ net1279 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ net1806 net538 net599 _05876_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12305_ net1304 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13285_ net1332 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
X_10497_ net134 net1027 net903 net1689 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15024_ clknet_leaf_61_wb_clk_i _02744_ _01389_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12236_ net1666 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08910__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net1630 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10552__A2 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ net829 _06557_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__and2_2
XANTENNA__09307__A _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _06795_ net479 net445 net1809 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a22o_1
X_15182__1563 vssd1 vssd1 vccd1 vccd1 _15182__1563/HI net1563 sky130_fd_sc_hd__conb_1
XFILLER_0_127_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11049_ net655 net706 _06527_ net824 vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__and4_1
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11275__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07705__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07181__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11572__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14808_ clknet_leaf_61_wb_clk_i net1830 _01173_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11291__B _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14412__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14739_ clknet_leaf_122_wb_clk_i _02503_ _01104_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10188__A _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08260_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07211_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\] net737
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__o221a_1
XANTENNA__13499__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ net1208 _04131_ _04132_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11511__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11568__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07142_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__or3_1
XANTENNA__14562__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07641__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07073_ _03011_ _03014_ net815 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10791__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11740__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\]
+ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or2_1
XANTENNA__08121__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09714_ _05073_ _05586_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__a21bo_1
X_06926_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\]
+ net876 _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07960__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ _05552_ _05586_ net580 vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__mux2_2
X_06857_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__and4b_4
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1292_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ net582 _05504_ _05505_ _05516_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11256__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08527_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\]
+ net971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout815_A _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08458_ net867 _04396_ _04399_ _04393_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08672__A1 net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _03341_ _03350_ net718 _03333_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_19_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08389_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[121\] net927
+ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10420_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _06139_ vssd1 vssd1
+ vccd1 vccd1 _06242_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09621__B1 _05562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ team_03_WB.instance_to_wrap.core.pc.current_pc\[24\] _06185_ net676 vssd1
+ vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13070_ net1285 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10282_ _03313_ _05972_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XANTENNA__08730__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08188__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net615 _06582_ net457 net365 net2301 vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__a32o_1
XANTENNA__07935__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A _05068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07573__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _03064_ vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout571 _03024_ vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
Xfanout582 net583 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_4
Xfanout593 net594 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_4
X_13972_ clknet_leaf_90_wb_clk_i _01736_ _00337_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12923_ net1361 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12039__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ net1344 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11805_ net2654 _06631_ net333 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12785_ net1315 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14524_ clknet_leaf_128_wb_clk_i _02288_ _00889_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ net593 net265 net477 _06808_ net1853 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a32o_1
XANTENNA__08905__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07871__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14455_ clknet_leaf_74_wb_clk_i _02219_ _00820_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ net2707 _06519_ net349 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XANTENNA__11331__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ net1402 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XANTENNA__08415__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10618_ net2325 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] net836 vssd1 vssd1 vccd1
+ vccd1 _02510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08415__B2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14386_ clknet_leaf_105_wb_clk_i _02150_ _00751_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11598_ net297 net2464 net454 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10549_ net1134 team_03_WB.instance_to_wrap.core.d_hit _02837_ vssd1 vssd1 vccd1
+ vccd1 _06292_ sky130_fd_sc_hd__nor3_4
XFILLER_0_109_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13337_ net1284 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11970__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ net1324 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15007_ clknet_leaf_39_wb_clk_i net55 _01372_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11567__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12219_ net1791 vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13199_ net1388 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07077__S1 net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11722__A1 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__C net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\]
+ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07691_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\] net758
+ net1037 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__o21a_1
X_09430_ net554 _04863_ _05042_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11506__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13802__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ _05294_ _05298_ _05293_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__o21a_1
XANTENNA__11238__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11789__A1 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08312_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\] net925
+ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09292_ _04893_ _05219_ _05215_ _04953_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13952__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\]
+ net946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\] net929
+ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__o221a_1
XANTENNA__10068__D team_03_WB.instance_to_wrap.core.decoder.inst\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08174_ net1057 _04112_ _04115_ net1201 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08116__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__and3_1
XANTENNA__11410__A0 _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1040_A _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11961__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07056_ _02996_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XANTENNA__12072__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11908__C _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XANTENNA__10516__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1305_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A1 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XANTENNA__11196__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ net723 _03899_ _03883_ _03882_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__o2bb2a_4
X_06909_ net1186 net883 vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07889_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[207\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\] net732
+ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10819__A3 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout932_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11416__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08342__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09628_ _05102_ _05104_ net565 vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a21o_1
XANTENNA__11643__C net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11229__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ _05302_ _05305_ _05187_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12570_ net1370 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
XANTENNA__07448__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08952__C _04893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11521_ _06381_ net649 _06634_ _06394_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__or4b_4
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14240_ clknet_leaf_133_wb_clk_i _02004_ _00605_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[594\]
+ sky130_fd_sc_hd__dfrtp_1
X_11452_ net650 _06577_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
X_15181__1562 vssd1 vssd1 vccd1 vccd1 _15181__1562/HI net1562 sky130_fd_sc_hd__conb_1
XFILLER_0_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10403_ _06227_ _06228_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] net678
+ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11401__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10204__A1 _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14171_ clknet_leaf_34_wb_clk_i _01935_ _00536_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09070__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ net712 _06527_ net697 vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__and3_1
XANTENNA__12771__A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__A1 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ net282 _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__nand2_1
XANTENNA_input61_A gpio_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ net1349 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08460__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13053_ net1375 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
X_10265_ _06089_ _06103_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_30_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1300 net1302 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__buf_4
X_12004_ net263 _06756_ net470 net450 net2189 vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__a32o_1
Xfanout1311 net1316 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1322 net1323 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__buf_4
X_10196_ net589 net659 vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1333 net1334 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07384__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1344 net1345 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__buf_4
XANTENNA__11180__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1355 net1358 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__buf_4
Xfanout1366 net1367 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13825__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08696__A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1377 net1380 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__buf_4
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_4
Xfanout1388 net1391 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__buf_4
Xfanout1399 net1405 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__buf_4
XFILLER_0_92_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13955_ clknet_leaf_19_wb_clk_i _01719_ _00320_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07136__A1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06928__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12906_ net1257 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
XANTENNA__13107__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13886_ clknet_leaf_48_wb_clk_i _01650_ _00251_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12837_ net1274 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08636__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12768_ net1378 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
X_14507_ clknet_leaf_36_wb_clk_i _02271_ _00872_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ net2173 net302 net342 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__mux2_1
XANTENNA__11640__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12699_ net1365 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ clknet_leaf_79_wb_clk_i _02202_ _00803_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput43 gpio_in[18] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11996__S net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput54 gpio_in[29] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
Xhold805 team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\] vssd1
+ vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
Xinput65 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14369_ clknet_leaf_0_wb_clk_i _02133_ _00734_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput76 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold816 team_03_WB.instance_to_wrap.core.register_file.registers_state\[332\] vssd1
+ vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11943__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput98 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
Xhold827 team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\] vssd1
+ vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07775__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 team_03_WB.instance_to_wrap.core.register_file.registers_state\[829\] vssd1
+ vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\] vssd1
+ vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11297__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08930_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\] net1204
+ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09364__A2 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\] net1075
+ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a221o_1
XANTENNA__07375__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _03749_ _03753_ _03752_ net1110 vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__a2bb2o_1
X_08792_ net921 _04732_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ net1083 net888 team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\]
+ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07127__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__B2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13017__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__o221a_1
XFILLER_0_79_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09413_ net576 _04832_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__nor2_1
XANTENNA__07015__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1088_A _02787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08627__A1 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _03170_ _03989_ _05149_ net606 vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a31o_1
XANTENNA__08545__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06854__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09230__A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11631__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ _04954_ _05215_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12067__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08226_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\]
+ net973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\] net1212
+ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__o221a_1
XANTENNA__10095__B _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ net1220 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\]
+ net949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__o221a_1
XANTENNA__09052__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1422_A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\] net746
+ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__a221oi_1
X_08088_ net1145 net1017 net682 vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07039_ net809 _02979_ _02980_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10050_ net6 net1032 net906 net2804 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o22a_1
XANTENNA__08012__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__S1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13998__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__B2 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_5_wb_clk_i _01504_ _00105_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08410__S0 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ net686 _05768_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11870__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ clknet_leaf_69_wb_clk_i _01435_ _00036_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10883_ net831 _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__nor2_4
XFILLER_0_109_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08079__C1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ net1340 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XANTENNA__08618__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11622__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12553_ net1252 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08094__A2 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10976__A2 _05142_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11504_ _06622_ net2684 net396 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ net1298 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ clknet_leaf_98_wb_clk_i _01987_ _00588_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ net1240 _06449_ net649 net701 vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__or4_4
XFILLER_0_106_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07595__A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11366_ net518 net641 _06735_ net408 net2151 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14154_ clknet_leaf_3_wb_clk_i _01918_ _00519_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ net1314 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
X_10317_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06152_ vssd1 vssd1
+ vccd1 vccd1 _06158_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ net714 _06557_ net825 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__and3_1
X_14085_ clknet_leaf_108_wb_clk_i _01849_ _00450_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ _04294_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] net670 vssd1
+ vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13036_ net1303 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XANTENNA__11689__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11153__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1130 net1133 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1141 team_03_WB.instance_to_wrap.core.decoder.inst\[23\] vssd1 vssd1 vccd1
+ vccd1 net1141 sky130_fd_sc_hd__buf_8
X_10179_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__inv_2
Xfanout1152 net1155 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_8
Xfanout1163 net1198 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
Xfanout1174 net1177 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10900__A2 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1185 net1197 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09315__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1196 net1197 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
XANTENNA__07761__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07109__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14987_ clknet_leaf_107_wb_clk_i net35 _01352_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ clknet_leaf_102_wb_clk_i _01702_ _00303_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11283__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09969__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13869_ clknet_leaf_104_wb_clk_i _01633_ _00234_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15108__1489 vssd1 vssd1 vccd1 vccd1 _15108__1489/HI net1489 sky130_fd_sc_hd__conb_1
X_07390_ _03328_ _03329_ _03330_ _03331_ net815 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08609__A1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11613__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[687\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[655\] net1006 net941
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08490__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\]
+ net771 net1122 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09034__A1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10924__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold602 team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\] vssd1
+ vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold613 team_03_WB.instance_to_wrap.CPU_DAT_I\[28\] vssd1 vssd1 vccd1 vccd1 net2197
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold624 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\] vssd1
+ vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08242__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold635 team_03_WB.instance_to_wrap.core.register_file.registers_state\[259\] vssd1
+ vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold646 team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\] vssd1
+ vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11392__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\] vssd1
+ vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold668 net128 vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09962_ _05885_ net1741 net292 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold679 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\] vssd1
+ vssd1 vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08913_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\]
+ net959 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09893_ _04031_ _04323_ net541 vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07348__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ net861 _04784_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__and3_1
XANTENNA__07443__S1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15180__1561 vssd1 vssd1 vccd1 vccd1 _15180__1561/HI net1561 sky130_fd_sc_hd__conb_1
X_08775_ _04715_ _04716_ net854 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout463_A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _03665_ _03667_ net1154 vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11852__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ net1130 _03589_ _03593_ _03596_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout630_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1372_A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout728_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07588_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\]
+ net881 vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10818__B _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10407__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11604__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ _05265_ _05267_ _05249_ _05253_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07284__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09258_ _03866_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\]
+ net955 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux2_1
X_09189_ net441 net433 _04565_ net548 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11907__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _06456_ _06503_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__nor2_1
XANTENNA__07036__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08784__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ net495 net646 _06652_ net417 net1838 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10102_ _05925_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11082_ net827 net301 vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__and2_2
XFILLER_0_120_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07339__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ clknet_leaf_38_wb_clk_i _00004_ _01275_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10033_ net25 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1
+ vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XANTENNA__09135__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ clknet_leaf_55_wb_clk_i _02605_ _01206_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12096__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14772_ clknet_leaf_61_wb_clk_i _02536_ _01137_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11984_ net301 net2727 net448 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__mux2_1
X_13723_ clknet_leaf_29_wb_clk_i _01487_ _00088_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11843__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10935_ net315 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[7\]
+ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__o31a_1
XANTENNA__07511__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11604__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ clknet_leaf_83_wb_clk_i _01418_ _00019_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10866_ net495 _06454_ net594 net521 net2097 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a32o_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ net1381 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13585_ net1282 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ net688 _05429_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07275__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12536_ net1362 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08913__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12467_ net1261 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_14206_ clknet_leaf_50_wb_clk_i _01970_ _00571_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ net299 net2682 net402 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__mux2_1
XANTENNA__09567__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12020__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15186_ net1567 vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_2
X_12398_ net1338 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11374__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08775__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14137_ clknet_leaf_103_wb_clk_i _01901_ _00502_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\]
+ sky130_fd_sc_hd__dfrtp_1
X_11349_ net1243 net833 net302 net667 vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__and4_1
XFILLER_0_123_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ clknet_leaf_91_wb_clk_i _01832_ _00433_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08527__B1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ net1361 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
X_06890_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _02832_ sky130_fd_sc_hd__nand2_2
XFILLER_0_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ net867 _04496_ _04501_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10637__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_07511_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\]
+ net879 _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a31o_1
X_08491_ net942 _04431_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__o21a_1
XANTENNA__14669__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11514__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07442_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[500\] net1144
+ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ net1090 net894 team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\]
+ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08689__S0 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13693__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ net1058 _05052_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07266__B1 _03207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11062__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08463__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09043_ net439 net431 _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\] vssd1
+ vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12011__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14049__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 team_03_WB.instance_to_wrap.CPU_DAT_I\[19\] vssd1 vssd1 vccd1 vccd1 net2005
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07569__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold432 team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\] vssd1
+ vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\] vssd1
+ vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _02601_ vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold465 team_03_WB.instance_to_wrap.core.register_file.registers_state\[441\] vssd1
+ vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11188__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold476 team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\] vssd1
+ vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 _02611_ vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1218_A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold498 team_03_WB.instance_to_wrap.core.register_file.registers_state\[230\] vssd1
+ vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 _02844_ vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09945_ _03425_ net660 vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__nor2_1
Xfanout912 net257 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09881__C _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 net924 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_4
XANTENNA_fanout580_A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 net936 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout678_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 _04087_ vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14199__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__buf_4
X_09876_ net542 _05816_ net664 vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a21bo_1
Xhold1110 team_03_WB.instance_to_wrap.core.register_file.registers_state\[599\] vssd1
+ vssd1 vccd1 vccd1 net2694 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout978 net979 vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_2
Xfanout989 net992 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\] vssd1
+ vssd1 vccd1 vccd1 net2705 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1132 team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\] vssd1
+ vssd1 vccd1 vccd1 net2716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08827_ team_03_WB.instance_to_wrap.core.decoder.inst\[18\] _04761_ net843 vssd1
+ vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a21o_1
Xhold1143 team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\] vssd1
+ vssd1 vccd1 vccd1 net2727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout845_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\] vssd1
+ vssd1 vccd1 vccd1 net2738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[704\] vssd1
+ vssd1 vccd1 vccd1 net2749 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07741__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\] vssd1
+ vssd1 vccd1 vccd1 net2760 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[333\] vssd1
+ vssd1 vccd1 vccd1 net2771 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08758_ net1214 _04698_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__and3_1
Xhold1198 team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\] vssd1
+ vssd1 vccd1 vccd1 net2782 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ net807 _03646_ _03647_ _03650_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08689_ _04627_ _04628_ _04629_ _04630_ net860 net922 vssd1 vssd1 vccd1 vccd1 _04631_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10720_ net528 _06350_ _06351_ net533 net2247 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07203__A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09246__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10651_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] team_03_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ net841 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ net1905 net536 net597 _03488_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a22o_1
X_13370_ net1324 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08454__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ net1290 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15040_ clknet_leaf_54_wb_clk_i _02760_ _01405_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09549__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12002__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ net1355 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08757__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net303 net2613 net493 vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12183_ net1662 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10564__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07655__S1 _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net1039 net832 net278 net666 vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__and4_1
X_15107__1488 vssd1 vssd1 vccd1 vccd1 _15107__1488/HI net1488 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11395__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11065_ _06609_ net2323 net423 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ net98 net97 net69 net68 vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14811__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12069__A0 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14824_ clknet_leaf_56_wb_clk_i net1954 _01189_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10619__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11816__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14755_ clknet_leaf_122_wb_clk_i net1711 _01120_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11842__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ net638 _06744_ net478 net371 net2438 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__B2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11292__A1 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13706_ clknet_leaf_9_wb_clk_i _01470_ _00071_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10918_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[10\] net307 vssd1
+ vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__nand2_1
XANTENNA__07496__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ clknet_leaf_42_wb_clk_i _02450_ _01051_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net640 _06707_ net480 net379 net1964 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__a32o_1
XANTENNA__11831__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07113__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13637_ net1421 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10849_ _06394_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07248__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08445__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ net1331 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08996__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12519_ net1398 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10474__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13499_ net1323 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11289__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15169_ net1550 vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11898__A3 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07783__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07991_ _02872_ _03931_ _03932_ _02870_ _03930_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__o221a_1
XANTENNA__13909__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _05669_ _05670_ net578 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06942_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\]
+ net773 vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09173__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09661_ net577 _05527_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__o21ai_1
X_06873_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ _02807_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__or3_1
XFILLER_0_119_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08612_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\]
+ net973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\] net938
+ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09592_ net577 _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09503__A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[638\] net1067
+ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08474_ _04080_ _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11822__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07023__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ _03364_ _03366_ net1151 vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11190__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1070_A net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__C _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[732\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\] net738
+ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1276_A team_03_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07287_ _03226_ _03228_ net809 vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1335_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ net1062 _04965_ _04966_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11338__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\] vssd1
+ vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold251 team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\] vssd1
+ vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _02633_ vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11889__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 net187 vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold284 net206 vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold295 team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\] vssd1
+ vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout962_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07962__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 _02863_ vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11419__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 net735 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_4
X_09928_ _05868_ net1917 net292 vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
Xfanout742 net751 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_4
Xfanout753 net755 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_2
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__clkbuf_4
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
Xfanout786 net787 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__buf_4
X_09859_ _05730_ _05746_ _05800_ _05757_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__or4b_1
XFILLER_0_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11365__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__S1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07175__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12870_ net1416 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11821_ net647 _06651_ net458 net328 net1824 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07478__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14540_ clknet_leaf_7_wb_clk_i _02304_ _00905_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\]
+ sky130_fd_sc_hd__dfrtp_1
X_11752_ _06576_ net468 net339 net2688 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a22o_1
XANTENNA__11381__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11813__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10703_ net525 _06339_ _06340_ net530 team_03_WB.instance_to_wrap.ADR_I\[27\] vssd1
+ vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a32o_1
XFILLER_0_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14471_ clknet_leaf_64_wb_clk_i _02235_ _00836_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11683_ _06725_ net391 net346 net2049 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ net1393 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XANTENNA_input91_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net1914 net842 vssd1
+ vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11026__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13353_ net1279 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
X_10565_ net1841 net536 net597 _05875_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ net1417 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07650__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13284_ net1392 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10496_ net104 net1027 net902 net1608 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a22o_1
X_15023_ clknet_leaf_33_wb_clk_i _02743_ _01388_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11131__C_N net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ net1617 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10537__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ net1642 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11329__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ _06632_ net2450 net422 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12097_ _06794_ net476 net445 net1866 vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11048_ net2554 net426 _06601_ net517 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07705__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09170__A3 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14807_ clknet_leaf_62_wb_clk_i net1816 _01172_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11572__B net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ net1390 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11291__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ clknet_leaf_120_wb_clk_i _02502_ _01103_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08666__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11999__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14669_ clknet_leaf_106_wb_clk_i _02433_ _01034_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12684__A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07210_ _03146_ _03151_ net816 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__mux2_1
XANTENNA__08418__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14707__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08190_ net1055 _04129_ _04130_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08969__B1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ net1189 net879 team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a21o_1
XANTENNA__11568__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09091__C1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07072_ net808 _03012_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10528__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11740__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\]
+ net897 _03915_ net1127 vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o311a_1
XANTENNA__13881__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09932__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ _05551_ _05654_ _05653_ _05652_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__o211a_1
X_06925_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\]
+ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout376_A _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__A3 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _04269_ _04326_ _04448_ _04386_ net556 net568 vssd1 vssd1 vccd1 vccd1 _05586_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06856_ net1414 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ net582 _05504_ _05505_ _05516_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__a31oi_2
XANTENNA__10379__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11256__A1 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ net859 _04464_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10059__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08657__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_A net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ net1055 _04397_ _04398_ net1201 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15106__1487 vssd1 vssd1 vccd1 vccd1 _15106__1487/HI net1487 sky130_fd_sc_hd__conb_1
XANTENNA_fanout808_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07408_ net718 _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08283__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ net942 _04328_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07339_ net1078 net885 team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\]
+ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__o21a_1
XANTENNA__09621__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _06184_ _06183_ net282 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09009_ net867 _04949_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or3b_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _05975_ _06111_ _06120_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__a31o_1
XANTENNA__10519__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08188__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12020_ net615 _06581_ net457 net365 net2358 vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__a32o_1
XANTENNA__07935__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A2 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout550 net552 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout572 net575 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
Xfanout583 _02950_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__buf_4
X_13971_ clknet_leaf_111_wb_clk_i _01735_ _00336_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__B2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _06464_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
XANTENNA__07699__A0 _03638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ net1372 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__09152__A3 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12853_ net1262 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ net2664 net264 net333 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12784_ net1428 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14523_ clknet_leaf_30_wb_clk_i _02287_ _00888_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11735_ net1902 net296 net342 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07598__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14454_ clknet_leaf_93_wb_clk_i _02218_ _00819_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07871__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11666_ net2373 _06628_ net350 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__mux2_1
X_13405_ net1326 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
X_10617_ net1654 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] net837 vssd1 vssd1 vccd1
+ vccd1 _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14385_ clknet_leaf_97_wb_clk_i _02149_ _00750_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11597_ net270 net2703 net452 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__mux2_1
X_13336_ net1291 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10548_ _06287_ _06290_ _06291_ team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1
+ vccd1 _02567_ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ net1259 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
X_10479_ net2717 net1026 net902 team_03_WB.instance_to_wrap.ADR_I\[27\] vssd1 vssd1
+ vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15006_ clknet_leaf_125_wb_clk_i net54 _01371_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_12218_ net1613 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11567__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ net1281 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11722__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__C_N _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net1638 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09128__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A3 _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07690_ _03630_ _03631_ net1152 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07272__S net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11238__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _05278_ _05281_ _05301_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08639__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08892__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\]
+ net985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\] net944
+ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__o221a_1
XANTENNA__09300__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09291_ _05227_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__nand2_1
XANTENNA__07311__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08654__A2 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08242_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\]
+ net946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[114\] net913
+ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__o221a_1
XANTENNA__07862__B1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09064__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\] net1209
+ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07614__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ net611 _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__A1 net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\] net1122
+ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a221o_1
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_113_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1033_A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XANTENNA__09228__A _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XANTENNA_fanout493_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XANTENNA__11196__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10921__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08590__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ net1111 _03897_ _03898_ _03894_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout660_A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ net1103 net899 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nor2_1
XANTENNA__10601__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\]
+ net880 _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__a31o_1
XANTENNA__08342__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09627_ net576 _05568_ _05566_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__o21ai_1
X_06839_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1 vccd1 vccd1
+ _02782_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout925_A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _05479_ _05499_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08509_ net937 _04449_ _04450_ net854 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09489_ _05332_ _05430_ _05324_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _06633_ net2542 net396 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07849__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11451_ net2710 net398 _06764_ net499 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10402_ net285 _06142_ _06224_ net678 vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__o31a_1
XFILLER_0_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10204__A2 _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ clknet_leaf_19_wb_clk_i _01934_ _00535_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\]
+ sky130_fd_sc_hd__dfrtp_1
X_11382_ net513 net639 _06743_ net407 net2198 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ net1266 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XANTENNA__07081__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10333_ _06118_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07357__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input54_A gpio_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13052_ net1350 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
X_10264_ _06092_ _06102_ _06104_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11704__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _06541_ net2337 net451 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__mux2_1
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__buf_4
Xfanout1312 net1316 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__buf_4
X_10195_ _06035_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1323 net1328 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__buf_4
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1334 net1335 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__buf_4
Xfanout1345 net1359 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__buf_2
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1356 net1357 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1367 net1387 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__clkbuf_2
Xfanout380 _06813_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1378 net1380 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__buf_4
Xfanout1389 net1390 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__buf_4
Xfanout391 net392 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_4
XANTENNA__11607__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ clknet_leaf_129_wb_clk_i _01718_ _00319_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14552__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09530__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ net1253 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
X_13885_ clknet_leaf_67_wb_clk_i _01649_ _00250_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12836_ net1306 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08916__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08097__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10979__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ net1374 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
XANTENNA__09833__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14506_ clknet_leaf_3_wb_clk_i _02270_ _00871_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11718_ net2016 _06434_ net342 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__mux2_1
X_15149__1530 vssd1 vssd1 vccd1 vccd1 _15149__1530/HI net1530 sky130_fd_sc_hd__conb_1
X_12698_ net1370 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14437_ clknet_leaf_123_wb_clk_i _02201_ _00802_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\]
+ sky130_fd_sc_hd__dfrtp_1
X_11649_ net2503 _06615_ net348 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__mux2_1
XANTENNA__09046__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12962__A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput44 gpio_in[19] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 gpio_in[30] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
X_14368_ clknet_leaf_133_wb_clk_i _02132_ _00733_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput66 wb_rst_i vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_1
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold806 team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\] vssd1
+ vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xinput77 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_2
Xhold817 team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\] vssd1
+ vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ net1326 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
Xhold828 team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\] vssd1
+ vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09698__A1_N _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput99 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_1
Xhold839 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\] vssd1
+ vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ clknet_leaf_27_wb_clk_i _02063_ _00664_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11297__B _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14082__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08860_ net1053 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\]
+ net1007 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\] net1207
+ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08572__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07375__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15105__1486 vssd1 vssd1 vccd1 vccd1 _15105__1486/HI net1486 sky130_fd_sc_hd__conb_1
X_07811_ net1123 _03751_ net1156 vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\] net998 net938
+ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o221a_1
XANTENNA__11517__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07742_ net1083 _02795_ net888 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__or3_1
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11459__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A0 _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08324__B2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\] net1115
+ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__o221a_1
XANTENNA__08875__A2 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09412_ _05350_ _05353_ _03025_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ _05283_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07835__B1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _04953_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07669__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08225_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[817\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\]
+ net973 vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1150_A team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ net1220 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\] net1066
+ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06870__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07107_ _03046_ _03048_ net1110 _03044_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ net721 _03999_ _04007_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__o31a_2
XFILLER_0_43_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1415_A net1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07038_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[227\] net730
+ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11147__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout875_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08012__B1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _04927_ _04930_ net863 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07771__C1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08315__A1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07118__A2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[4\] net308 net684 vssd1
+ vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__a21o_1
XANTENNA__08410__S1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ clknet_leaf_74_wb_clk_i _01434_ _00035_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10882_ net690 _06475_ _06476_ _06474_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__a31o_2
XFILLER_0_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12621_ net1301 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09815__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12552_ net1352 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XANTENNA__07826__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11503_ _06479_ net2612 net394 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12483_ net1300 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14222_ clknet_leaf_69_wb_clk_i _01986_ _00587_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\]
+ sky130_fd_sc_hd__dfrtp_1
X_11434_ net266 net2626 net404 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__mux2_1
XANTENNA__11386__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07054__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ clknet_leaf_59_wb_clk_i _01917_ _00518_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\]
+ sky130_fd_sc_hd__dfrtp_1
X_11365_ net1244 net834 net300 net667 vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ net1427 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
X_10316_ net282 _06128_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and3_1
X_14084_ clknet_leaf_15_wb_clk_i _01848_ _00449_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11296_ net511 net637 _06715_ net415 net2259 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13035_ net1275 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
X_10247_ _05986_ _05991_ _06086_ _05988_ _05983_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__o311ai_4
XFILLER_0_119_37 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1120 _02785_ vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08554__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1131 net1133 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09751__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1142 net1144 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
X_10178_ _03242_ _06018_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__and3_1
XANTENNA__10361__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1153 net1155 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_4
XANTENNA__13942__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_2
Xfanout1175 net1177 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1186 net1187 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_2
XANTENNA__09729__S1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
X_14986_ clknet_leaf_123_wb_clk_i net65 _01351_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12102__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13937_ clknet_leaf_94_wb_clk_i _01701_ _00302_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13868_ clknet_leaf_5_wb_clk_i _01632_ _00233_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12819_ net1265 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13799_ clknet_leaf_69_wb_clk_i _01563_ _00164_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07817__A0 _03756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09282__A2 _05146_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ net1129 _03950_ _03951_ net1111 _03949_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__a311o_1
XANTENNA__11800__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10924__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold603 team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\] vssd1
+ vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07045__A1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold614 team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\] vssd1
+ vssd1 vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\] vssd1
+ vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\] vssd1
+ vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\] vssd1
+ vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08793__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold658 team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\] vssd1
+ vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09961_ _03678_ net660 vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold669 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\] vssd1
+ vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08912_ net1199 _04850_ _04853_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__or3_1
XFILLER_0_102_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09892_ _05182_ _05502_ _05503_ net591 vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__a211o_1
X_08843_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[224\] net927
+ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10888__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07899__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10151__S net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08774_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\]
+ net974 team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\] net938
+ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09940__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[653\]
+ net727 _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout456_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07505__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07656_ net1107 _03597_ net1130 vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06865__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout623_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _03526_ _03528_ net608 vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15195__1573 vssd1 vssd1 vccd1 vccd1 _15195__1573/HI net1573 sky130_fd_sc_hd__conb_1
XFILLER_0_113_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1365_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09326_ _05265_ _05267_ _05253_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09895__B _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ _04072_ _05147_ net606 vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08481__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08208_ _04120_ _04149_ net551 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09188_ _05128_ _05129_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11368__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout992_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ net1077 net1012 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net703 _06468_ net695 vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__and3_1
XANTENNA__10591__A1 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13965__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _05921_ _05922_ _05941_ _05944_ _05920_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a221o_4
X_11081_ _06618_ net2350 net423 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07339__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10032_ net26 net1032 net906 net2692 vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__o22a_1
XANTENNA__11540__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ clknet_leaf_55_wb_clk_i net2081 _01205_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09135__B _05076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ clknet_leaf_62_wb_clk_i _02535_ _01136_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11983_ net302 net2839 net450 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__mux2_1
XANTENNA__08839__A2 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08395__S0 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ clknet_leaf_22_wb_clk_i _01486_ _00087_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_10934_ net686 _05730_ _06399_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13653_ clknet_leaf_89_wb_clk_i _01417_ _00018_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10865_ net653 net705 _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12604_ net1347 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13584_ net1278 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10796_ net281 net2737 net522 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ net1413 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
XANTENNA__07275__A1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104__1485 vssd1 vssd1 vccd1 vccd1 _15104__1485/HI net1485 sky130_fd_sc_hd__conb_1
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14740__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ net1410 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14205_ clknet_leaf_76_wb_clk_i _01969_ _00570_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\]
+ sky130_fd_sc_hd__dfrtp_1
X_11417_ net271 net2490 net401 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__mux2_1
XANTENNA__12020__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15185_ net1566 vssd1 vssd1 vccd1 vccd1 la_data_out[121] sky130_fd_sc_hd__buf_2
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12397_ net1291 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14136_ clknet_leaf_12_wb_clk_i _01900_ _00501_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11348_ net515 net635 _06726_ net408 net2074 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a32o_1
XANTENNA__10582__B2 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14067_ clknet_leaf_111_wb_clk_i _01831_ _00432_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10760__A _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ net713 _06513_ net825 vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__and3_1
XANTENNA__08527__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13018_ net1366 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XANTENNA__09724__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11531__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11067__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14969_ clknet_leaf_33_wb_clk_i _02721_ _01334_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07510_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\]
+ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08490_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\] net988 net928
+ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a221o_1
XANTENNA__08376__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07441_ net1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[372\] net1116
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07372_ _03312_ _03313_ net608 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11598__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08689__S1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ net1212 _05050_ _05051_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__and3_1
XANTENNA__07266__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11062__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ net843 _04970_ _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08405__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold400 team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\] vssd1
+ vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12011__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold411 team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\] vssd1
+ vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _02590_ vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07569__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08766__A1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 net156 vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 net233 vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold455 team_03_WB.instance_to_wrap.core.register_file.registers_state\[634\] vssd1
+ vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11188__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold466 team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\] vssd1
+ vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 net174 vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__B2 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07974__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout902 net904 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_2
X_09944_ _05876_ net2133 net295 vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
Xhold488 team_03_WB.instance_to_wrap.CPU_DAT_I\[27\] vssd1 vssd1 vccd1 vccd1 net2072
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10670__A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout913 net915 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_4
Xhold499 team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\] vssd1
+ vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1113_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 _04088_ vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout946 net948 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout957 net968 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08140__A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _03604_ _04820_ _05069_ _03601_ net1018 vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__a32o_1
Xhold1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\] vssd1
+ vssd1 vccd1 vccd1 net2684 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 _04086_ vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_2
Xhold1111 team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\] vssd1
+ vssd1 vccd1 vccd1 net2695 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout979 net980 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_4
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08826_ net1214 _04763_ _04764_ _04767_ net1077 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 team_03_WB.instance_to_wrap.core.register_file.registers_state\[142\] vssd1
+ vssd1 vccd1 vccd1 net2706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 net122 vssd1 vssd1 vccd1 vccd1 net2717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15128__1509 vssd1 vssd1 vccd1 vccd1 _15128__1509/HI net1509 sky130_fd_sc_hd__conb_1
Xhold1144 team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\] vssd1
+ vssd1 vccd1 vccd1 net2728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\] vssd1
+ vssd1 vccd1 vccd1 net2739 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07741__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\] vssd1
+ vssd1 vccd1 vccd1 net2750 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[739\] net923
+ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a221o_1
Xhold1177 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\] vssd1
+ vssd1 vccd1 vccd1 net2761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\] vssd1
+ vssd1 vccd1 vccd1 net2772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1199 team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\] vssd1
+ vssd1 vccd1 vccd1 net2783 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ net739 _03648_ _03649_ net802 vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11825__A1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08688_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__mux2_1
XANTENNA__07190__S net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\]
+ net873 _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11006__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] team_03_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ net841 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11589__A0 _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09309_ _02938_ _05126_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__nor2_1
X_10581_ net2036 net536 net597 _03458_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12320_ net1408 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XANTENNA__13221__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12002__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ net1362 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11379__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A0 _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__A0 _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08757__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ net279 net2640 net490 vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__mux2_1
X_12182_ net1744 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11761__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net2154 net420 _06642_ net515 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
XANTENNA__11676__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08509__A1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11395__B net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ net1240 _06449_ net628 _06463_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__or4_2
XFILLER_0_60_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ net78 net67 net92 net89 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08390__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07732__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14823_ clknet_leaf_55_wb_clk_i net1781 _01188_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08196__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14754_ clknet_leaf_119_wb_clk_i _02518_ _01119_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11966_ net638 _06743_ net479 net372 net2298 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13705_ clknet_leaf_77_wb_clk_i _01469_ _00070_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ net692 _05686_ net587 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07496__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14685_ clknet_leaf_42_wb_clk_i _02449_ _01050_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11292__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ net624 _06706_ net459 net377 net2674 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ net1329 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10848_ _06381_ _06390_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09920__C_N _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ net1404 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10779_ net1039 _02808_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07799__A2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08996__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12518_ net1419 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13498_ net1326 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12449_ net1290 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XANTENNA__11289__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15168_ net1549 vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11752__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__C1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14119_ clknet_leaf_64_wb_clk_i _01883_ _00484_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07783__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\]
+ net784 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15099_ net1480 vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_2
XANTENNA__07420__B2 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06941_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[900\]
+ net773 vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__mux2_1
XANTENNA__11504__A0 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09660_ net577 _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__nand2_1
X_06872_ _02811_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\] net998
+ net921 _04552_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ _05393_ _05418_ net570 vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13660__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13306__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\] net1202
+ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07304__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ net845 _04414_ _04401_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10491__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\]
+ net886 _03365_ net1144 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07239__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[636\] net724
+ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__o221a_1
XFILLER_0_128_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout321_A net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07286_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[137\] net778
+ net733 _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a211o_1
XANTENNA__11991__A0 _06487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\]
+ net982 net1071 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12880__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1230_A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1328_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__A0 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold230 net189 vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\] vssd1
+ vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[25\] vssd1 vssd1 vccd1
+ vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\] vssd1
+ vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout788_A net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold274 team_03_WB.instance_to_wrap.CPU_DAT_I\[21\] vssd1 vssd1 vccd1 vccd1 net1858
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\] vssd1
+ vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold296 team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\] vssd1
+ vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout710 net711 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
Xfanout721 _02863_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07962__A2 _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout732 net734 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_09927_ _03638_ net660 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout743 net745 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout955_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_2
Xfanout776 net785 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09858_ _05768_ _05784_ _05798_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__or3_1
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__buf_4
X_15103__1484 vssd1 vssd1 vccd1 vccd1 _15103__1484/HI net1484 sky130_fd_sc_hd__conb_1
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__buf_4
XANTENNA__07175__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08911__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08372__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\]
+ net976 net1072 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__mux4_1
X_09789_ _05250_ _05269_ _05246_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11820_ net651 _06650_ net461 net328 net1856 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ _06574_ net473 net339 net2571 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
XANTENNA__11274__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ _06311_ _06337_ net600 vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10482__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14470_ clknet_leaf_79_wb_clk_i _02234_ _00835_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\]
+ sky130_fd_sc_hd__dfrtp_1
X_11682_ _06724_ net386 net344 net2730 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ net1309 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11026__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10633_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] team_03_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ net842 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14509__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13352_ net1284 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
X_10564_ net1951 net535 net596 _05874_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a22o_1
XANTENNA_input84_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11982__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12303_ net1377 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
X_13283_ net1392 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ net105 net1027 net902 net1881 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ clknet_leaf_55_wb_clk_i _02742_ _01387_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dfrtp_1
X_12234_ net1691 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07884__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11734__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12165_ net1679 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07953__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net829 net267 vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__and2_2
X_12096_ _06793_ net482 net446 net2102 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a22o_1
XANTENNA__09155__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13683__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ net642 _06600_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08363__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09604__A _05545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06913__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13126__A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14806_ clknet_leaf_39_wb_clk_i _02570_ _01171_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11572__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12998_ net1411 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737_ clknet_leaf_117_wb_clk_i _02501_ _01102_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08666__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ net640 _06726_ net480 net371 net1957 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14668_ clknet_leaf_5_wb_clk_i _02432_ _01033_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\]
+ sky130_fd_sc_hd__dfstp_1
X_13619_ net1329 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
XANTENNA__08418__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14189__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14599_ clknet_leaf_64_wb_clk_i _02363_ _00964_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15127__1508 vssd1 vssd1 vccd1 vccd1 _15127__1508/HI net1508 sky130_fd_sc_hd__conb_1
XFILLER_0_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11973__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[226\] net735
+ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07641__B2 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10932__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11725__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11740__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07973_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\]
+ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09146__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ net584 _04775_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__or2_2
XFILLER_0_103_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06924_ net1098 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\]
+ net1148 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07157__B1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09643_ _05185_ _05501_ _05192_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06855_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[29\] vssd1 vssd1 vccd1
+ vccd1 _02798_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout369_A net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ net359 _05508_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08525_ net854 _04465_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__or3_1
XANTENNA__07034__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11256__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08657__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout536_A net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1180_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10464__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07969__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[860\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\] net1208
+ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__o221a_1
XANTENNA__08564__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07407_ net1140 _03347_ _03348_ net1157 _03346_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o311a_1
XANTENNA__07880__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ net1238 team_03_WB.instance_to_wrap.core.register_file.registers_state\[185\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[153\] net990 net927
+ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07338_ _03277_ _03279_ net608 vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__mux2_2
XFILLER_0_89_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11964__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14801__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07632__A1 net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[969\]
+ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ net915 _04947_ _04948_ net856 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10280_ _03822_ _06117_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11731__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _04821_ vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_4
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
Xfanout562 _03063_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
X_13970_ clknet_leaf_103_wb_clk_i _01734_ _00335_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout573 net575 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07148__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout584 _02892_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
Xfanout595 net599 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_4
X_12921_ net1355 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08896__B1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12852_ net1322 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net2583 _06630_ net335 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12783_ net1377 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
XANTENNA__12785__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08982__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11734_ net593 _06519_ net476 _06808_ net1849 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a32o_1
X_14522_ clknet_leaf_6_wb_clk_i _02286_ _00887_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07320__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07871__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ net2218 _06627_ net348 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__mux2_1
X_14453_ clknet_leaf_87_wb_clk_i _02217_ _00818_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13404_ net1324 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
X_10616_ net1715 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] net837 vssd1 vssd1 vccd1
+ vccd1 _02512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14384_ clknet_leaf_82_wb_clk_i _02148_ _00749_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\]
+ sky130_fd_sc_hd__dfrtp_1
X_11596_ _06504_ net2333 net454 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11955__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14481__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ net1285 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
X_10547_ team_03_WB.instance_to_wrap.wb.curr_state\[0\] _06284_ _06289_ vssd1 vssd1
+ vccd1 vccd1 _06291_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13266_ net1422 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XANTENNA__11970__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10478_ net123 net1026 net904 net1736 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08503__A _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15005_ clknet_leaf_125_wb_clk_i net53 _01370_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_12217_ net1733 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
X_13197_ net1320 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
XANTENNA__11567__C net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__B1 _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11183__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ net1643 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11722__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12079_ net625 _06643_ net463 net447 net1852 vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__B1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08639__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08892__B net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08310_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\] net983
+ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__or2_1
XANTENNA__11803__S net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A1 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__nand2_1
XANTENNA__07311__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ net929 _04181_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__o21a_1
XANTENNA__11104__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08172_ net1055 _04111_ _04113_ net1066 vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__a211o_1
XANTENNA__09064__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102__1483 vssd1 vssd1 vccd1 vccd1 _15102__1483/HI net1483 sky130_fd_sc_hd__conb_1
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11946__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07123_ net1178 net1013 _02835_ net1246 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07614__A1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07054_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\] net1146
+ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11961__A3 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_28_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XANTENNA__11477__C _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__B _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XANTENNA__07917__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XANTENNA__11196__D net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout486_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ net728 _03886_ _03887_ net1140 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a211o_1
XANTENNA__09244__A _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06907_ net1158 net879 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__nand2_8
X_07887_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[79\]
+ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout653_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ net573 _05483_ _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__a21oi_2
X_06838_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[8\] vssd1 vssd1 vccd1
+ vccd1 _02781_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09557_ net591 _05430_ _05480_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__o31a_2
XANTENNA_fanout820_A _02846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08508_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[671\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\] net920
+ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _05306_ _05307_ _05311_ _05329_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o31a_1
XFILLER_0_52_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10988__B2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08439_ net863 _04380_ _04375_ net846 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ net628 _06575_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__and2_1
XANTENNA__11937__A0 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ net285 _06226_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__S0 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08802__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ net712 net296 net698 vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ net1411 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
X_10332_ _05975_ _06111_ _06116_ _06114_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__a31o_1
XANTENNA__11952__A3 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09419__A _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ net1361 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10263_ _06097_ _06100_ _06096_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__C _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12002_ net264 _06756_ net475 net451 net2118 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a32o_1
Xfanout1302 net1317 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__buf_2
XANTENNA__08030__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _04565_ net673 _06033_ _02893_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o211a_1
XANTENNA_input47_A gpio_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1313 net1314 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__buf_4
Xfanout1324 net1328 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__buf_4
Xfanout1335 net1433 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__buf_2
Xfanout1346 net1349 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__buf_4
Xfanout1357 net1358 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__buf_4
Xfanout370 _06815_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_4
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1368 net1373 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__buf_4
Xfanout381 net384 vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_6
Xfanout1379 net1380 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__buf_2
Xfanout392 _06802_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__clkbuf_8
X_13953_ clknet_leaf_2_wb_clk_i _01717_ _00318_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15126__1507 vssd1 vssd1 vccd1 vccd1 _15126__1507/HI net1507 sky130_fd_sc_hd__conb_1
XFILLER_0_96_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09530__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ net1286 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ clknet_leaf_119_wb_clk_i _01648_ _00249_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08993__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ net1296 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08097__A1 net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12766_ net1383 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14505_ clknet_leaf_59_wb_clk_i _02269_ _00870_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07402__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ net1970 net276 net342 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__mux2_1
XANTENNA__11640__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ net1358 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11648_ net2600 _06614_ net349 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__mux2_1
XANTENNA__09046__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14436_ clknet_leaf_16_wb_clk_i _02200_ _00801_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
XFILLER_0_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09597__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 gpio_in[0] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput45 gpio_in[20] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10763__A _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ clknet_leaf_109_wb_clk_i _02131_ _00732_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[721\]
+ sky130_fd_sc_hd__dfrtp_1
X_11579_ _06418_ net2741 net452 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
Xinput56 gpio_in[31] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xhold807 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\] vssd1
+ vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput78 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput89 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
X_13318_ net1284 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
Xhold818 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\] vssd1
+ vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11943__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold829 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\] vssd1
+ vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
X_14298_ clknet_leaf_19_wb_clk_i _02062_ _00663_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07775__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14227__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11297__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ net1265 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__B2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07810_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[427\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[299\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\]
+ net770 net1121 vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__mux4_1
X_08790_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[546\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\]
+ net974 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12105__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08309__C1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__B1 _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ net1170 net874 _02796_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11459__A2 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07672_ net806 _03609_ _03610_ _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _05351_ _05352_ net556 vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07015__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ _04207_ _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__nand2_1
XANTENNA__08088__A1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11092__A0 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07835__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ _03790_ _05214_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11631__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09938__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08224_ net1059 _04165_ _04164_ net1070 vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _04097_ sky130_fd_sc_hd__nand2_4
XANTENNA_fanout401_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10198__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1143_A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07106_ net1156 _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08086_ net1139 _04017_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[67\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[99\] net746
+ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1310_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08012__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout770_A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout868_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10612__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08988_ net856 _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and3_1
X_07939_ net1121 _03877_ _03878_ net1111 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10658__A0 team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10950_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[4\] net306 vssd1 vssd1
+ vccd1 vccd1 _06533_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09609_ net574 _04535_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__nand2_2
X_10881_ net690 _06475_ _06476_ _06474_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input101_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ net1298 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
XANTENNA__08079__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09276__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__A2 _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ net1398 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XANTENNA__11622__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11502_ _06621_ net2759 net393 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__mux2_1
X_12482_ net1365 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09123__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ net267 net2831 net403 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__mux2_1
X_14221_ clknet_leaf_105_wb_clk_i _01985_ _00586_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11386__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ clknet_leaf_27_wb_clk_i _01916_ _00517_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\]
+ sky130_fd_sc_hd__dfrtp_1
X_11364_ net515 net634 _06734_ net408 net2139 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__a32o_1
XANTENNA__11398__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10315_ _05969_ _06127_ _05970_ _05964_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__a211o_1
X_13103_ net1391 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14083_ clknet_leaf_19_wb_clk_i _01847_ _00448_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ net715 _06550_ net824 vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__and3_1
XANTENNA__08988__A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13034_ net1258 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
X_10246_ _05987_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nor2_1
XANTENNA__11689__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1110 net1111 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__buf_4
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
XANTENNA__09751__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__C_N net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1132 net1133 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_4
XANTENNA__07211__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _04922_ net673 vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__or2_1
XANTENNA__08199__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 net1155 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10361__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_2
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__clkbuf_2
Xfanout1187 net1196 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_2
X_14985_ clknet_leaf_107_wb_clk_i net64 _01350_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1198 team_03_WB.instance_to_wrap.core.decoder.inst\[20\] vssd1 vssd1 vccd1
+ vccd1 net1198 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15101__1482 vssd1 vssd1 vccd1 vccd1 _15101__1482/HI net1482 sky130_fd_sc_hd__conb_1
X_13936_ clknet_leaf_82_wb_clk_i _01700_ _00301_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[290\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08711__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13867_ clknet_leaf_18_wb_clk_i _01631_ _00232_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12818_ net1412 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13798_ clknet_leaf_74_wb_clk_i _01562_ _00163_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07817__A1 _03758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11613__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ net1301 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09019__B1 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10821__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__B2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09114__S0 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ clknet_leaf_115_wb_clk_i _02183_ _00784_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[773\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10924__C net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07278__S net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08242__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold604 team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\] vssd1
+ vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold615 team_03_WB.instance_to_wrap.core.register_file.registers_state\[44\] vssd1
+ vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\] vssd1
+ vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold637 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\] vssd1
+ vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\] vssd1
+ vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09960_ _05884_ net1767 net294 vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__mux2_1
Xhold659 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\] vssd1
+ vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08911_ net935 _04852_ _04851_ net1056 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__o211a_1
XFILLER_0_102_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09891_ _05825_ _05826_ _05832_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07202__C1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08842_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\] net943
+ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__a221o_1
XANTENNA__09742__B2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08773_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\] net999
+ net921 _04714_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07724_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[685\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__B1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07655_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[942\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[814\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[782\]
+ net760 _02785_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10668__A _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout351_A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1093_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07586_ net682 _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__and2b_1
XFILLER_0_53_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08138__A _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11065__A0 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09325_ _05253_ _05266_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout616_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10812__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1358_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _05196_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07284__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__C net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08207_ net438 net436 _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nor3_2
XFILLER_0_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09187_ net441 net433 _04592_ net553 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__o31a_1
XFILLER_0_7_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10607__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ _04075_ net436 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__or2_2
XANTENNA__11907__A3 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125__1506 vssd1 vssd1 vccd1 vccd1 _15125__1506/HI net1506 sky130_fd_sc_hd__conb_1
XFILLER_0_71_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08233__A1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07441__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ net727 _04008_ _04009_ net1108 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__a31o_1
XANTENNA__07992__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10100_ _02831_ _02926_ _05940_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__o31a_1
XFILLER_0_124_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11080_ net830 net302 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and2_2
XFILLER_0_41_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10031_ team_03_WB.instance_to_wrap.BUSY_O net1036 team_03_WB.instance_to_wrap.wb.prev_BUSY_O
+ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__or3b_4
XFILLER_0_105_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13219__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11540__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08941__C1 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ clknet_leaf_38_wb_clk_i _02534_ _01135_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.WRITE_I
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12096__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ net275 net2743 net450 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08395__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ clknet_leaf_84_wb_clk_i _01485_ _00086_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ net512 net593 _06519_ net522 net1876 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07511__A3 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13652_ clknet_leaf_91_wb_clk_i _01416_ _00017_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10864_ net1246 _02808_ net1245 vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__or3b_4
XFILLER_0_131_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14072__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ net1364 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13583_ net1282 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
X_10795_ net684 _06398_ net586 _06402_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__o211a_2
XANTENNA__12793__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07887__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10803__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12534_ net1341 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07680__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ net1304 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14204_ clknet_leaf_128_wb_clk_i _01968_ _00569_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[558\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11416_ net300 net2342 net404 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__mux2_1
XANTENNA__08224__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09421__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12396_ net1300 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
X_15184_ net1565 vssd1 vssd1 vccd1 vccd1 la_data_out[120] sky130_fd_sc_hd__buf_2
XFILLER_0_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11347_ net275 net713 net698 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__and3_1
X_14135_ clknet_leaf_74_wb_clk_i _01899_ _00500_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14066_ clknet_leaf_101_wb_clk_i _01830_ _00431_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\]
+ sky130_fd_sc_hd__dfrtp_1
X_11278_ net497 net620 _06706_ net413 net2361 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a32o_1
XANTENNA__09724__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] net670 vssd1 vssd1 vccd1
+ vccd1 _06071_ sky130_fd_sc_hd__nand2_1
XANTENNA__13129__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ net1357 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07735__B1 _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 team_03_WB.instance_to_wrap.SEL_I\[0\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14968_ clknet_leaf_32_wb_clk_i _02720_ _01333_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09342__A _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ clknet_leaf_116_wb_clk_i _01683_ _00284_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[273\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11834__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ clknet_leaf_37_wb_clk_i _02662_ _01264_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11083__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07440_ _03378_ _03381_ net816 vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net1017 net682 vssd1
+ vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09110_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[430\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\]
+ net955 net1069 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14565__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08463__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__A2 _03205_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09041_ net864 _04981_ _04982_ net847 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_894 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08215__A1 _04084_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\] vssd1
+ vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__A2 _06569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold412 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\] vssd1
+ vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_03_WB.instance_to_wrap.core.register_file.registers_state\[314\] vssd1
+ vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _02599_ vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\] vssd1
+ vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold456 team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\] vssd1
+ vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10573__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 team_03_WB.instance_to_wrap.core.register_file.registers_state\[296\] vssd1
+ vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold478 team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\] vssd1
+ vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _04029_ net662 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold489 team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\] vssd1
+ vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 net927 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09715__A1 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout936 _04087_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_2
Xfanout947 net948 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
X_09874_ _03604_ _05069_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__nand2_1
XANTENNA__07726__B1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout958 net959 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__clkbuf_4
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1106_A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[483\] vssd1
+ vssd1 vccd1 vccd1 net2685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\] vssd1
+ vssd1 vccd1 vccd1 net2696 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ _04765_ _04766_ net1060 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a21o_1
Xhold1123 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\] vssd1
+ vssd1 vccd1 vccd1 net2707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 _02630_ vssd1 vssd1 vccd1 vccd1 net2718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\] vssd1
+ vssd1 vccd1 vccd1 net2729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout566_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1156 team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\] vssd1
+ vssd1 vccd1 vccd1 net2740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[516\] vssd1
+ vssd1 vccd1 vccd1 net2751 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12078__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\] vssd1
+ vssd1 vccd1 vccd1 net2762 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[579\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\] net939
+ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\] vssd1
+ vssd1 vccd1 vccd1 net2773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10089__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07707_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\]
+ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__or2_1
XANTENNA__11286__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__A2 _06656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[808\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[776\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout733_A net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07638_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\]
+ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ net1187 net883 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\]
+ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11721__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13502__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _04565_ _05248_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__nand2_1
X_10580_ net2032 net535 net596 _05890_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
XANTENNA__08454__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10845__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07500__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09239_ _05180_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12118__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11022__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ net1371 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__inv_2
X_15100__1481 vssd1 vssd1 vccd1 vccd1 _15100__1481/HI net1481 sky130_fd_sc_hd__conb_1
XANTENNA__12002__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _06413_ net2729 net491 vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__mux2_1
XANTENNA__11210__A0 _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12181_ net1597 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10564__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A1 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ net634 _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__A _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\] vssd1
+ vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ net830 net281 vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__and2_2
XFILLER_0_25_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11395__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ net94 net93 net96 net95 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07193__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08390__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__B2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822_ clknet_leaf_57_wb_clk_i _02586_ _01187_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14753_ clknet_leaf_128_wb_clk_i _02517_ _01118_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11816__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ net636 _06742_ net476 net371 net1950 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ clknet_leaf_18_wb_clk_i _01468_ _00069_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14588__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ net506 net593 _06505_ net522 net1935 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14684_ clknet_leaf_42_wb_clk_i _02448_ _01049_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08693__A1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11896_ net639 _06705_ net476 net379 net2445 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13635_ net1313 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10847_ net274 net2489 net524 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08445__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07248__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ net1400 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ net1245 net1246 net1015 vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_67_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__C1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12517_ net1275 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08540__S1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ net1323 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12448_ net1413 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11289__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11201__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ net1548 vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_2
X_12379_ net1362 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ clknet_leaf_77_wb_clk_i _01882_ _00483_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15098_ net1479 vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_2
XFILLER_0_10_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06940_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\]
+ net773 vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14049_ clknet_leaf_2_wb_clk_i _01813_ _00414_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07708__B1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06871_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nand4_4
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11806__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08610_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\] net973
+ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or2_1
X_09590_ _05420_ _05525_ net570 vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11268__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ net1208 _04482_ _04481_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15124__1505 vssd1 vssd1 vccd1 vccd1 _15124__1505/HI net1505 sky130_fd_sc_hd__conb_1
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11107__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08472_ _04408_ _04413_ net867 vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07423_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\]
+ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or2_1
XANTENNA__09800__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07023__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07354_ _03294_ _03295_ net812 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07285_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[169\]
+ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08135__B _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1056_A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09946__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 net106 vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 team_03_WB.instance_to_wrap.CPU_DAT_I\[0\] vssd1 vssd1 vccd1 vccd1 net1815
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10681__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\] vssd1
+ vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold253 net176 vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09247__A _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\] vssd1
+ vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _02592_ vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 net203 vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout700 _06561_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_8
Xhold297 team_03_WB.instance_to_wrap.ADR_I\[11\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout711 _06460_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_2
X_09926_ _05861_ net1940 net293 vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_8
Xfanout733 net734 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 net745 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__clkbuf_4
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_2
Xfanout766 net767 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_2
X_09857_ _05784_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__or2_1
Xfanout777 net779 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07175__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout788 net800 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
Xfanout799 net800 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_2
XANTENNA_fanout948_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08372__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08808_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a221o_1
XANTENNA__10620__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ net583 _05720_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a21oi_4
X_08739_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\] net975
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08124__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11017__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _06573_ net482 net338 net2363 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
XANTENNA__07478__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10701_ _06316_ _06338_ net604 vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11681_ _06723_ net390 net346 net2021 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ net1313 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08427__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10632_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] team_03_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ net842 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11431__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13351_ net1330 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
X_10563_ net1777 net535 net596 _05873_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12302_ net1336 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ net1804 net1025 net902 team_03_WB.instance_to_wrap.ADR_I\[12\] vssd1 vssd1
+ vccd1 vccd1 _02615_ sky130_fd_sc_hd__a22o_1
X_13282_ net1392 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07650__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input77_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15021_ clknet_leaf_61_wb_clk_i _02741_ _01386_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12233_ net1747 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08286__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10537__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11734__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12164_ net1653 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10942__C1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ net263 net2394 net423 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ net620 _06666_ net459 net444 net1986 vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09591__S net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ net702 net714 net296 vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__or3b_1
XFILLER_0_99_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14805_ clknet_leaf_56_wb_clk_i _02569_ _01170_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11572__D net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ net1277 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14736_ clknet_leaf_122_wb_clk_i _02500_ _01101_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07124__B _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ net643 _06725_ net483 net371 net2088 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08666__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14667_ clknet_leaf_38_wb_clk_i _02431_ _01032_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11879_ net617 _06688_ net456 net377 net2120 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a32o_1
X_13618_ net1402 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XANTENNA__08418__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ clknet_leaf_79_wb_clk_i _02362_ _00963_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07140__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11422__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13549_ net1307 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
XANTENNA__09091__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12981__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11973__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07070_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[98\] net745
+ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a221o_1
XFILLER_0_67_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08670__S net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14603__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15219_ net911 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10528__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11725__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07972_ net808 _03909_ _03910_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o22a_1
X_09711_ _03682_ net540 _05041_ _03679_ _02804_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__o32a_1
XANTENNA__11489__A0 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06923_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\]
+ net876 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07157__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09642_ _05185_ _05192_ _05501_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__and3_1
XANTENNA__13317__A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ net1 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__inv_2
XANTENNA__10161__B1 _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06857__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09573_ net326 _05354_ _05384_ _05513_ _05512_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08524_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\]
+ net971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[255\] net937
+ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__o221a_1
XANTENNA__08657__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09854__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[828\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[796\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1173_A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06873__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout529_A _02923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07406_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\] net1146
+ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08386_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[25\]
+ net990 vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1281_A team_03_WB.instance_to_wrap.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07337_ team_03_WB.instance_to_wrap.core.decoder.inst\[29\] net1016 net682 vssd1
+ vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11964__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07985__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07268_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\]
+ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or2_1
XANTENNA__11003__C net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout898_A net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ _04945_ _04946_ net850 vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07199_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\]
+ net753 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__mux2_1
XANTENNA__10615__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10519__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A1 _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 net533 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_4
X_09909_ _05454_ _05563_ _05848_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or4_1
XANTENNA__09705__A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout552 _03105_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09910__C_N _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07148__A1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout585 _02891_ vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
Xfanout596 net598 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
X_12920_ net1369 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12851_ net1259 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ net2276 net265 net333 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12782_ net1336 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14521_ clknet_leaf_103_wb_clk_i _02285_ _00886_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07856__C1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ net2163 net297 net342 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ clknet_leaf_92_wb_clk_i _02216_ _00817_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\]
+ sky130_fd_sc_hd__dfrtp_1
X_11664_ net2416 _06505_ net349 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08056__A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13403_ net1402 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07608__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10615_ net1681 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] net836 vssd1 vssd1 vccd1
+ vccd1 _02513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ clknet_leaf_97_wb_clk_i _02147_ _00748_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\]
+ sky130_fd_sc_hd__dfrtp_1
X_11595_ _06499_ net2659 net453 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13334_ net1318 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10546_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265_ net1315 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10477_ net124 net1026 net902 net1633 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123__1504 vssd1 vssd1 vccd1 vccd1 _15123__1504/HI net1504 sky130_fd_sc_hd__conb_1
X_15004_ clknet_leaf_124_wb_clk_i net52 _01369_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_12216_ net1768 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ net1299 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XANTENNA__11567__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11183__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12147_ net1693 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07119__B _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__B1 net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12078_ _06783_ net480 net446 net1963 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a22o_1
X_11029_ net701 net709 net299 vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07135__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__A net1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08639__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14719_ clknet_leaf_123_wb_clk_i _02483_ _01084_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08240_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\] net946 net913
+ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11104__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\]
+ net949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\] net1209
+ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__o221a_1
XANTENNA__09064__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08498__S0 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11946__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09496__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ net611 _03059_ _03061_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08811__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10943__B _06527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10084__A_N _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07053_ net611 _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07090__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_11_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11120__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08024__C1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XANTENNA__07378__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__D _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XANTENNA__11174__A2 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1019_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ net1117 _03896_ _03895_ net1130 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout381_A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06868__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06906_ net1114 net895 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07886_ net732 _03824_ _03825_ _03826_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a32o_1
X_09625_ net567 net557 _05137_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__and3_1
XANTENNA__11882__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 _02780_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout646_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1388_A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _05371_ _05485_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06884__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[575\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__mux2_1
XANTENNA__14649__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11634__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout813_A _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _05389_ _05390_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a21o_2
XFILLER_0_77_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10988__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08438_ _04376_ _04377_ _04379_ _04378_ net933 net857 vssd1 vssd1 vccd1 vccd1 _04380_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09055__A1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\] net935
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13673__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14799__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ _06076_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07066__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ net512 net636 _06742_ net407 net1757 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ team_03_WB.instance_to_wrap.core.pc.current_pc\[27\] _06150_ vssd1 vssd1
+ vccd1 vccd1 _06169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_666 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11030__A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ _05981_ _06091_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__nand2_1
XANTENNA__14029__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13050_ net1366 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07369__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11387__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _06532_ net2783 net450 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__mux2_1
X_10193_ _06033_ _06034_ _02893_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__a21oi_1
Xfanout1303 net1305 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__buf_4
Xfanout1314 net1315 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__buf_4
Xfanout1325 net1328 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__buf_2
Xfanout1336 net1337 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__buf_4
Xfanout1347 net1349 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__buf_2
XANTENNA__08318__B1 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1358 net1359 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__buf_2
Xfanout360 _04776_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1369 net1373 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__buf_4
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13952_ clknet_leaf_130_wb_clk_i _01716_ _00317_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout393 net394 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_6
X_12903_ net1399 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11873__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ clknet_leaf_25_wb_clk_i _01647_ _00248_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07541__A1 net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ net1364 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08485__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09818__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10428__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11625__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12765_ net1370 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14504_ clknet_leaf_34_wb_clk_i _02268_ _00869_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\]
+ sky130_fd_sc_hd__dfrtp_1
X_11716_ net2280 _06426_ net341 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12696_ net1371 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14435_ clknet_leaf_26_wb_clk_i _02199_ _00800_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09046__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11647_ net2773 _06613_ net348 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14366_ clknet_leaf_48_wb_clk_i _02130_ _00731_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[720\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput35 gpio_in[10] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
X_11578_ _06413_ net2719 net452 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__mux2_1
Xinput46 gpio_in[21] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10763__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput57 gpio_in[32] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold808 team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\] vssd1
+ vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10600__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13317_ net1294 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
X_10529_ net137 net1023 net1019 net1774 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
Xinput79 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_1
Xhold819 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\] vssd1
+ vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14297_ clknet_leaf_112_wb_clk_i _02061_ _00662_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13248_ net1410 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11156__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ net1360 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XANTENNA__08021__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07765__D1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11086__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07740_ _03680_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__or2_2
XANTENNA__07207__S1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire614_A _02842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11864__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ net738 _03611_ _03612_ net801 vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__a31o_1
X_09410_ net546 _04149_ _04209_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09809__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11616__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _04207_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07296__B1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08493__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09272_ _03244_ _05145_ net607 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14941__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_115_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08223_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\]
+ net973 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10954__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12041__A0 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__A2 _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ team_03_WB.instance_to_wrap.core.decoder.inst\[19\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _04096_ sky130_fd_sc_hd__and2_1
XANTENNA__08424__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06870__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[481\]
+ net876 _03045_ net1125 vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__a311o_1
X_08085_ net1133 _04022_ _04024_ _04026_ net721 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__o41a_1
XFILLER_0_114_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11488__C net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07036_ _02975_ _02977_ net803 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout596_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__A2 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08548__B1 net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14321__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__B1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\] net914
+ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a221o_1
XANTENNA__07771__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ net1157 _03879_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11855__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07869_ net1113 _03809_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11724__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _05464_ _05470_ net571 vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ net315 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\]
+ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__or4b_1
X_15122__1503 vssd1 vssd1 vccd1 vccd1 _15122__1503/HI net1503 sky130_fd_sc_hd__conb_1
XANTENNA__11607__A0 _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09539_ net581 _04824_ _05125_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12550_ net1419 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07287__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _06469_ net2825 net393 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10830__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[24\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12481_ net1290 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XANTENNA__10864__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14220_ clknet_leaf_7_wb_clk_i _01984_ _00585_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09123__S1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ net509 net263 _06756_ net403 net2191 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a32o_1
XANTENNA__12032__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07134__S0 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11386__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08787__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ clknet_leaf_65_wb_clk_i _01915_ _00516_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11363_ net716 net272 net699 vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13102_ net1337 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
X_10314_ _02766_ net675 _06133_ _06155_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14082_ clknet_leaf_129_wb_clk_i _01846_ _00447_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\]
+ sky130_fd_sc_hd__dfrtp_1
X_11294_ net509 net632 _06714_ net416 net2297 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ net1255 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10245_ _05991_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nor2_1
XANTENNA__09200__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08634__S0 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1100 net1105 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1111 net1114 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_8
X_10176_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] net673 vssd1 vssd1 vccd1
+ vccd1 _06018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1122 net1129 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_4
Xfanout1133 _02784_ vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_6
Xfanout1144 net1145 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_4
Xfanout1155 net1160 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1166 net1198 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_2
XANTENNA__12099__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_2
X_14984_ clknet_leaf_124_wb_clk_i net63 _01349_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1188 net1191 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_2
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11846__A0 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10649__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13935_ clknet_leaf_101_wb_clk_i _01699_ _00300_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__B1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07514__B2 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13866_ clknet_leaf_4_wb_clk_i _01630_ _00231_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12817_ net1312 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
X_13797_ clknet_leaf_107_wb_clk_i _01561_ _00162_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12748_ net1296 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12679_ net1398 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14418_ clknet_leaf_101_wb_clk_i _02182_ _00783_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12023__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08227__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08244__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14349_ clknet_leaf_106_wb_clk_i _02113_ _00714_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold605 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\] vssd1
+ vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold616 team_03_WB.instance_to_wrap.core.register_file.registers_state\[281\] vssd1
+ vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap324 _05746_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_2
Xhold627 team_03_WB.instance_to_wrap.core.register_file.registers_state\[291\] vssd1
+ vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold638 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\] vssd1
+ vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap357 _04863_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold649 team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\] vssd1
+ vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08910_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09890_ net325 _05437_ _05770_ net360 _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a221o_2
XFILLER_0_81_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08841_ _04781_ _04782_ net853 vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08772_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\] net974
+ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07723_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\] net763
+ net741 _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__a211o_1
XANTENNA__11837__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06939__S0 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07654_ net1107 _03594_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__or3_1
XANTENNA__08419__A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net1016 vssd1 vssd1 vccd1
+ vccd1 _03527_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1086_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09324_ net589 _05252_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09255_ _05069_ _05195_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nor2_1
XANTENNA__10684__A _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout511_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13060__A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout609_A _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _04134_ _04147_ net845 vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__mux2_8
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_133_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12014__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09186_ net441 net433 _04620_ net548 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08154__A team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08137_ _03567_ _04076_ _04077_ _04078_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_86_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1420_A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09430__A1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07441__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11011__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[726\]
+ net766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[758\] net740
+ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout880_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14837__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07992__A1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11719__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ _02959_ _02960_ net1110 vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10623__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ team_03_WB.instance_to_wrap.BUSY_O team_03_WB.instance_to_wrap.wb.prev_BUSY_O
+ net1034 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10879__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07744__A1 net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13861__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11828__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ net276 net2604 net450 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13235__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ clknet_leaf_12_wb_clk_i _01484_ _00085_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ net833 _06517_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__nor2_4
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14217__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ clknet_leaf_113_wb_clk_i _01415_ _00016_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10863_ net1246 _02809_ net1245 vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__and3b_1
XFILLER_0_131_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12602_ net1365 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13582_ net1281 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XANTENNA__11056__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ _05799_ _05867_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__A1 _02798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12533_ net1265 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12005__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12464_ net1417 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07680__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ clknet_leaf_28_wb_clk_i _01967_ _00568_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ net272 net2484 net404 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15183_ net1564 vssd1 vssd1 vccd1 vccd1 la_data_out[119] sky130_fd_sc_hd__buf_2
XANTENNA__10567__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ net1253 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12020__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ clknet_leaf_85_wb_clk_i _01898_ _00499_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_11346_ net519 net642 _06725_ net408 net2296 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07983__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ clknet_leaf_95_wb_clk_i _01829_ _00430_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09607__B _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08607__S0 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ net1242 net832 _06509_ net668 vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07408__A net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ net1369 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
X_10228_ _06004_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
XANTENNA__07735__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ _05041_ net659 vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__and2_1
Xhold2 team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\] vssd1
+ vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11819__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14967_ clknet_leaf_41_wb_clk_i _02719_ _01332_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13145__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13918_ clknet_leaf_58_wb_clk_i _01682_ _00283_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[272\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14898_ clknet_leaf_37_wb_clk_i _02661_ _01263_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08160__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13849_ clknet_leaf_93_wb_clk_i _01613_ _00214_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12984__A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__C1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ net720 _03311_ _03303_ _03296_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_70_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07120__C1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09040_ net870 _04973_ _04976_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__or3_1
XFILLER_0_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07671__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10558__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\] vssd1
+ vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 team_03_WB.instance_to_wrap.core.ru.state\[4\] vssd1 vssd1 vccd1 vccd1 net1997
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold424 team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\] vssd1
+ vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold435 team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\] vssd1
+ vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold446 team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\] vssd1
+ vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07974__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\] vssd1
+ vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold468 team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\] vssd1
+ vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__A2 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09942_ _05875_ net2425 net293 vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__mux2_1
X_15121__1502 vssd1 vssd1 vccd1 vccd1 _15121__1502/HI net1502 sky130_fd_sc_hd__conb_1
XFILLER_0_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold479 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\] vssd1
+ vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout904 _06285_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13884__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_2
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout926 net927 vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_4
Xfanout937 net945 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__clkbuf_4
X_09873_ net359 _05422_ _05814_ net585 vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__o22a_1
Xfanout948 net968 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08923__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
X_08824_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\]
+ net1001 team_03_WB.instance_to_wrap.core.register_file.registers_state\[737\] net1072
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a221o_1
Xhold1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\] vssd1
+ vssd1 vccd1 vccd1 net2686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\] vssd1
+ vssd1 vccd1 vccd1 net2697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1001_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\] vssd1
+ vssd1 vccd1 vccd1 net2708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\] vssd1
+ vssd1 vccd1 vccd1 net2719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_03_WB.instance_to_wrap.core.register_file.registers_state\[442\] vssd1
+ vssd1 vccd1 vccd1 net2730 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ net939 _04694_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
Xhold1157 team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\] vssd1
+ vssd1 vccd1 vccd1 net2741 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10679__A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout461_A net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\] vssd1
+ vssd1 vccd1 vccd1 net2752 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\] vssd1
+ vssd1 vccd1 vccd1 net2763 sky130_fd_sc_hd__dlygate4sd3_1
X_07706_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\]
+ net891 vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__or3_1
XANTENNA__11286__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08686_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\]
+ net978 vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__mux2_1
XANTENNA__11825__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07637_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\]
+ net1145 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1370_A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08439__C1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\] net798
+ net732 _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09100__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ _04565_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__nor2_1
XANTENNA__10618__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ _03433_ _03434_ _03439_ _03440_ net1111 net1131 vssd1 vssd1 vccd1 vccd1 _03441_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09238_ _04323_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11022__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ net441 net433 _04647_ net554 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__o31a_1
XFILLER_0_107_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12002__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ net280 net2620 net490 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA__07414__B1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ net1664 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07965__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ net713 net694 net303 vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 team_03_WB.instance_to_wrap.core.register_file.registers_state\[482\] vssd1
+ vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09167__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold991 team_03_WB.instance_to_wrap.core.register_file.registers_state\[705\] vssd1
+ vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ net2637 net427 _06608_ net519 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10013_ _03103_ net1868 net289 vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08390__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14821_ clknet_leaf_53_wb_clk_i net1771 _01186_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14752_ clknet_leaf_122_wb_clk_i _02516_ _01117_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11964_ net640 _06741_ net480 net371 net2111 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a32o_1
XANTENNA__08059__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13703_ clknet_leaf_69_wb_clk_i _01467_ _00068_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10915_ net833 _06503_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__nor2_2
X_14683_ clknet_leaf_53_wb_clk_i _02447_ _01048_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09890__A1 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11895_ net622 _06704_ net462 net377 net2196 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07350__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11912__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13634_ net1315 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10846_ _06443_ _06444_ _06445_ net587 vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13565_ net1402 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
X_10777_ net1246 net1015 vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nand2_2
XFILLER_0_125_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11213__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12516_ net1311 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07653__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ net1326 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ net1356 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07405__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ net1547 vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08602__C1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ net1372 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07956__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11752__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ clknet_leaf_108_wb_clk_i _01881_ _00482_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11329_ net263 net2627 net412 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__mux2_1
X_15097_ net1478 vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10960__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07138__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14048_ clknet_leaf_130_wb_clk_i _01812_ _00413_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07708__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09173__A3 _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[2\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08381__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07184__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11094__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11268__A1 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[798\]
+ net953 net1065 vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ net1208 _04411_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11107__B _06523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07304__C net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13603__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07422_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[884\]
+ net886 _03363_ net1116 vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__o311a_1
XANTENNA__07892__B1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07353_ net1106 _03291_ _03292_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09633__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07644__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07284_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[9\] net778
+ net749 _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09023_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\]
+ net982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\] net1071
+ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__o221a_1
XFILLER_0_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 team_03_WB.instance_to_wrap.ADR_I\[7\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 _02615_ vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 _02571_ vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold243 team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\] vssd1
+ vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\] vssd1
+ vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 team_03_WB.instance_to_wrap.core.register_file.registers_state\[392\] vssd1
+ vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_03_WB.instance_to_wrap.core.register_file.registers_state\[869\] vssd1
+ vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 team_03_WB.instance_to_wrap.CPU_DAT_I\[4\] vssd1 vssd1 vccd1 vccd1 net1871
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1216_A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10951__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09962__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout701 _06559_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_6
Xhold298 _02614_ vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _05646_ _05676_ _05856_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__and3_1
Xfanout712 net715 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_4
Xfanout723 _02863_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_8
XANTENNA__12889__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 net735 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout676_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 net751 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__clkbuf_4
Xfanout756 net760 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__clkbuf_4
Xfanout767 net785 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_2
X_09856_ _05080_ _05609_ _05791_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o211a_4
Xfanout778 net779 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10703__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 net800 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_4
XANTENNA__08372__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\] net1204
+ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__a221o_1
X_09787_ _02954_ _05508_ _05724_ _05728_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout843_A net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] _02832_ vssd1 vssd1 vccd1
+ vccd1 _02941_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08738_ net442 net434 net589 net547 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__o31a_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08669_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\]
+ net979 net1073 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11732__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ _02769_ _06315_ _02768_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10482__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ _06722_ net387 net344 net2025 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] team_03_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ net841 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11033__A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ net1277 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
X_10562_ net2134 net534 net595 _05872_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08832__C1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ net1318 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
X_13281_ net1392 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
X_10493_ net107 net1025 net905 net1789 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
X_15020_ clknet_leaf_62_wb_clk_i _02740_ _01385_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ net1749 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07884__C net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14405__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__C1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08286__S1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11734__A2 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12163_ net1645 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _06631_ net2800 net422 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12094_ _06792_ net470 net445 net1972 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12799__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09155__A3 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ net2763 net426 _06599_ net512 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a22o_1
XANTENNA__14555__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08363__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07166__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07797__S0 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06913__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14804_ clknet_leaf_39_wb_clk_i _02568_ _01169_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12996_ net1306 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08115__B2 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1091 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11947_ net625 _06724_ net463 net369 net2063 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32o_1
X_14735_ clknet_leaf_11_wb_clk_i _02499_ _01100_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11670__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ clknet_leaf_3_wb_clk_i _02430_ _01031_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ net625 _06687_ net464 net377 net2356 vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__a32o_1
X_15120__1501 vssd1 vssd1 vccd1 vccd1 _15120__1501/HI net1501 sky130_fd_sc_hd__conb_1
XFILLER_0_54_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07421__A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13617_ net1425 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10829_ net313 net311 net322 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__a31o_1
XANTENNA__09076__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14597_ clknet_leaf_124_wb_clk_i _02361_ _00962_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ net1325 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08823__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13479_ net1397 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15218_ net912 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14085__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11089__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07929__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__A2 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ net1530 vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10933__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07971_ net745 _03911_ _03912_ net805 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__a31o_1
X_09710_ _03682_ _05041_ _05651_ net664 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a22o_1
X_06922_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net873 vssd1 vssd1 vccd1
+ vccd1 _02864_ sky130_fd_sc_hd__nand2_8
XANTENNA__09000__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ net582 _05338_ _05564_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a31o_4
XFILLER_0_78_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06853_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[12\] vssd1
+ vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__inv_2
XANTENNA__13922__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11118__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09811__A net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ net1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[95\]
+ net971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\] net920
+ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__o221a_1
XANTENNA__07034__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11661__A1 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ net1055 _04394_ _04395_ net1065 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a211o_1
XANTENNA__07969__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07405_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[639\] net1122
+ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__o221a_1
X_08385_ _04150_ _04210_ _04269_ _04326_ net559 net568 vssd1 vssd1 vccd1 vccd1 _04327_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout424_A _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1166_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07617__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] net821 vssd1 vssd1 vccd1
+ vccd1 _03278_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07267_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11003__D net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07632__A3 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1333_A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09006_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\] net994 net931
+ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o221a_1
XANTENNA__09258__A _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07198_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\]
+ net752 vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout793_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09790__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _06448_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_4
Xfanout531 net533 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_2
XANTENNA__11727__S net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout542 _04815_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09908_ _05518_ _05583_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__nand3_1
XANTENNA__10631__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_2
Xfanout564 _03063_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
XANTENNA__08345__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout575 _03024_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_4
Xfanout597 net598 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__clkbuf_2
X_09839_ net580 _05778_ _05779_ _05780_ _05078_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a311o_1
XFILLER_0_57_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12850_ net1419 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net2263 _06629_ net333 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__mux2_1
XANTENNA__11101__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12781_ net1290 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XANTENNA__07305__C1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14520_ clknet_leaf_9_wb_clk_i _02284_ _00885_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11732_ net2372 net270 net341 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07320__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07241__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14451_ clknet_leaf_113_wb_clk_i _02215_ _00816_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09058__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11663_ net2311 _06626_ net348 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13402_ net1314 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10614_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\] net1823 net838
+ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__mux2_1
XANTENNA__07608__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ clknet_leaf_70_wb_clk_i _02146_ _00747_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11594_ net299 net2845 net453 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ net1321 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
X_10545_ team_03_WB.instance_to_wrap.wb.curr_state\[0\] _06288_ vssd1 vssd1 vccd1
+ vccd1 _06289_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ net1429 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10476_ net1845 net1026 net902 team_03_WB.instance_to_wrap.ADR_I\[30\] vssd1 vssd1
+ vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
XANTENNA__08072__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ clknet_leaf_123_wb_clk_i net51 _01368_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12215_ net1610 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__clkbuf_1
X_13195_ net1276 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07387__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12146_ net1637 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10391__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09128__A3 _05068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12077_ net618 _06640_ net460 net444 net2109 vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11028_ net499 net649 _06588_ net428 net2340 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a32o_1
XANTENNA__07416__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10143__A1 _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11891__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ net1259 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XANTENNA__10777__A net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13153__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14718_ clknet_leaf_39_wb_clk_i _02482_ _01083_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09049__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ clknet_leaf_104_wb_clk_i _02413_ _01014_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1003\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08170_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__mux2_1
XANTENNA__08681__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08498__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07121_ net611 _03059_ _03061_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08272__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09078__A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07052_ net1145 _02818_ net1015 net1039 vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08024__B1 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11120__B net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_100_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08575__A1 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_11_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08132__D _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13328__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[791\]
+ net785 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06868__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ net1141 net881 vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nand2_8
XANTENNA__06868__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\]
+ net880 net1149 vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout374_A _06814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07535__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ net576 _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__nand2_1
X_06836_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[17\] vssd1 vssd1 vccd1
+ vccd1 _02779_ sky130_fd_sc_hd__inv_2
XANTENNA__08856__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09555_ _04778_ _05106_ _05489_ _05492_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__o2111ai_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout541_A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__B team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1283_A net1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13063__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ net550 _04417_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__o21ai_2
XANTENNA__10880__D_N team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _05371_ _05404_ _05412_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14250__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout806_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08368_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\] net917
+ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07319_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\]
+ net874 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__and3_1
XANTENNA__10626__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08299_ _04239_ _04240_ net861 vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__B1 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10330_ team_03_WB.instance_to_wrap.core.pc.current_pc\[28\] _06168_ net675 vssd1
+ vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10261_ _06093_ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08566__A1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ net265 _06756_ net479 net451 net1981 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a32o_1
X_10192_ _04565_ net672 vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__or2_1
XANTENNA__08620__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1304 net1305 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__buf_4
Xfanout1315 net1316 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__buf_4
Xfanout1326 net1328 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__buf_4
Xfanout1337 net1339 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__buf_2
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08318__A1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1348 net1349 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__buf_4
Xfanout361 net362 vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_6
Xfanout1359 net1387 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__clkbuf_4
Xfanout372 _06815_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_8
Xfanout383 net384 vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_6
X_13951_ clknet_leaf_115_wb_clk_i _01715_ _00316_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[305\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout394 _06778_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07526__C1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ net1411 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13882_ clknet_leaf_21_wb_clk_i _01646_ _00247_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12833_ net1266 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11625__A1 _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12764_ net1350 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08067__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11715_ net2168 _06422_ net343 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__mux2_1
X_14503_ clknet_leaf_64_wb_clk_i _02267_ _00868_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12695_ net1415 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11920__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ net2453 _06612_ net348 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
X_14434_ clknet_leaf_128_wb_clk_i _02198_ _00799_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[788\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14743__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14365_ clknet_leaf_67_wb_clk_i _02129_ _00730_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08254__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput36 gpio_in[11] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ net280 net2591 net453 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 gpio_in[22] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 gpio_in[33] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10061__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13316_ net1294 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
Xinput69 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_1
X_10528_ net138 net1029 net1021 net1862 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold809 team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\] vssd1
+ vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
X_14296_ clknet_leaf_10_wb_clk_i _02060_ _00661_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13247_ net1376 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
X_10459_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] _06273_ net680 vssd1
+ vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11875__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ net1366 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XANTENNA__08530__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ net1618 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08309__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12105__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07670_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\]
+ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_1
XANTENNA__06985__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__A1 _02923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _03170_ _05151_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11040__C_N net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07296__A1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09271_ _05211_ _05212_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nand2_1
XANTENNA__08493__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08222_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\] net1213
+ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08705__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10954__B _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08153_ net855 _04091_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07048__B2 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11131__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__a221oi_1
XANTENNA__10052__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[790\] net789
+ net1037 _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11488__D _06463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07035_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\] net792
+ net731 _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1031_A _06283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1129_A _02785_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__A _05477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout491_A _06680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07756__C1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\] net931
+ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09970__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07937_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\]
+ net768 net1121 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux4_1
XANTENNA__14616__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08586__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[475\]
+ net781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[507\] net1149
+ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__o221a_1
XANTENNA__06895__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08720__A1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08181__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _05548_ _05371_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and2b_1
X_07799_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\] net796
+ net730 _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout923_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _05306_ _05307_ _05311_ _05329_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nor4_1
XFILLER_0_66_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10210__A _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08079__A3 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__A2 _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11025__B _06586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09469_ _05410_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11500_ _06454_ net2354 net393 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10830__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ net1408 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10864__B _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ net268 net2820 net403 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__S1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14150_ clknet_leaf_76_wb_clk_i _01914_ _00515_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ net500 net628 _06733_ net405 net1782 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ net1319 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ net283 _06154_ net675 vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ clknet_leaf_2_wb_clk_i _01845_ _00446_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14146__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ net1243 net834 _06545_ net669 vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13032_ net1351 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10244_ _05996_ _05999_ _06084_ _05994_ _05992_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__o311a_2
XANTENNA_input52_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11543__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08634__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1101 net1102 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_2
Xfanout1112 net1114 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ _03789_ _06015_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__xnor2_1
Xfanout1123 net1125 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__buf_4
Xfanout1134 _02765_ vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_4
Xfanout1145 team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1 vccd1
+ vccd1 net1145 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14296__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_4
Xfanout1167 net1168 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14983_ clknet_leaf_124_wb_clk_i net62 _01348_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1178 net1198 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
XANTENNA__11915__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1189 net1191 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
X_13934_ clknet_leaf_73_wb_clk_i _01698_ _00299_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08172__C1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08711__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ clknet_leaf_77_wb_clk_i _01629_ _00230_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ net1428 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13796_ clknet_leaf_12_wb_clk_i _01560_ _00161_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[150\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ net1254 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XANTENNA__11650__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12678_ net1419 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08525__A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09120__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11629_ _06703_ net386 net356 net2482 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a22o_1
XANTENNA__12023__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14417_ clknet_leaf_93_wb_clk_i _02181_ _00782_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09975__A0 _02921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__B1 _05907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08778__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14348_ clknet_leaf_8_wb_clk_i _02112_ _00713_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold606 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\] vssd1
+ vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10585__B2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 team_03_WB.instance_to_wrap.core.register_file.registers_state\[239\] vssd1
+ vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07450__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\] vssd1
+ vssd1 vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ clknet_leaf_65_wb_clk_i _02043_ _00644_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold639 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\] vssd1
+ vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09356__A _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08840_ net1236 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\]
+ net986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\] net941
+ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__o221a_1
XANTENNA__07202__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08771_ net553 _04712_ _04680_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07722_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and3_1
XANTENNA__11837__A1 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13663__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08702__A1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06939__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07653_ net1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\] net1117
+ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11126__A net1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07584_ net722 _03500_ _03506_ _03525_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o31a_4
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09323_ _05263_ _05264_ _05256_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10965__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout337_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1079_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _05069_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08205_ net863 _04145_ _04146_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09185_ _04824_ _04831_ _05126_ _05123_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a31o_1
XANTENNA__14169__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09966__A0 _05887_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1246_A team_03_WB.instance_to_wrap.core.decoder.inst\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _03352_ _03391_ _03428_ _03903_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__and4_1
XFILLER_0_114_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__B2 _05886_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07441__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08067_ net1171 team_03_WB.instance_to_wrap.core.register_file.registers_state\[598\]
+ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
XANTENNA__10904__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07018_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[899\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\]
+ net773 net1123 vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__mux4_1
XANTENNA__09266__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07729__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10879__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08941__A1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08969_ _04909_ _04910_ net1215 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11735__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ net278 net2801 net448 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10931_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11036__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13650_ clknet_leaf_100_wb_clk_i _01414_ _00015_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10862_ net1240 _06388_ _06459_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12601_ net1356 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
X_13581_ net1402 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XANTENNA__11056__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10793_ _05799_ _05867_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__and2b_2
XANTENNA__13251__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12532_ net1320 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12463_ net1410 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XANTENNA__07680__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11414_ net2494 net401 _06753_ net500 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14202_ clknet_leaf_20_wb_clk_i _01966_ _00567_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15182_ net1563 vssd1 vssd1 vccd1 vccd1 la_data_out[118] sky130_fd_sc_hd__buf_2
X_12394_ net1256 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
XANTENNA__09421__A2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07968__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ clknet_leaf_88_wb_clk_i _01897_ _00498_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\]
+ sky130_fd_sc_hd__dfrtp_1
X_11345_ net276 net714 net698 vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07395__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14064_ clknet_leaf_112_wb_clk_i _01828_ _00429_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11516__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ net510 net636 _06705_ net415 net2487 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a32o_1
XANTENNA__08607__S1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ net1416 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
X_10227_ _06009_ _06012_ _06065_ _06006_ _06002_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a311oi_2
XANTENNA__08393__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14931__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] net659 vssd1 vssd1 vccd1
+ vccd1 _06000_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold3 team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\] vssd1
+ vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11645__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14966_ clknet_leaf_56_wb_clk_i _02718_ _01331_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ net592 _05519_ _05540_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08145__C1 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13917_ clknet_leaf_60_wb_clk_i _01681_ _00282_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07043__S0 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14897_ clknet_leaf_37_wb_clk_i _02660_ _01262_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13848_ clknet_leaf_12_wb_clk_i _01612_ _00213_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08954__S net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08448__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13779_ clknet_leaf_113_wb_clk_i _01543_ _00144_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07120__B1 _03043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07671__A1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10007__A0 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10558__B2 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold403 team_03_WB.instance_to_wrap.CPU_DAT_I\[29\] vssd1 vssd1 vccd1 vccd1 net1987
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14461__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\] vssd1
+ vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold425 team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] vssd1 vssd1 vccd1 vccd1
+ net2009 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold436 team_03_WB.instance_to_wrap.core.register_file.registers_state\[187\] vssd1
+ vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold447 team_03_WB.instance_to_wrap.ADR_I\[19\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold458 team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\] vssd1
+ vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _03900_ net661 vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__nor2_1
Xhold469 team_03_WB.instance_to_wrap.core.register_file.registers_state\[761\] vssd1
+ vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11770__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10934__B1_N _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout905 _06285_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout916 _04088_ vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_4
Xfanout927 net928 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
X_09872_ _05734_ _05736_ net576 vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout938 net945 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__buf_4
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08823_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a221o_1
Xhold1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\] vssd1
+ vssd1 vccd1 vccd1 net2687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\] vssd1
+ vssd1 vccd1 vccd1 net2698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
Xhold1125 team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\] vssd1
+ vssd1 vccd1 vccd1 net2709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1136 team_03_WB.instance_to_wrap.core.register_file.registers_state\[143\] vssd1
+ vssd1 vccd1 vccd1 net2720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13336__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1147 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\] vssd1
+ vssd1 vccd1 vccd1 net2731 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[515\] net1001
+ net923 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__o21a_1
Xhold1158 team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\] vssd1
+ vssd1 vccd1 vccd1 net2742 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[731\] vssd1
+ vssd1 vccd1 vccd1 net2753 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\] net726
+ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__o221a_1
XANTENNA__11286__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[904\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout454_A net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07636_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\]
+ net873 vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__and3_1
XANTENNA__07053__B _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07567_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[568\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__or3_1
XANTENNA__10695__A _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1363_A net1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_A _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ net529 _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07498_ _03435_ _03436_ net746 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11994__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ _04032_ _05154_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07662__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07500__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11022__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ _05108_ _05109_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout990_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\]
+ net891 _04060_ net1143 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__o311a_1
XFILLER_0_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07414__A1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10634__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ net846 _05027_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__o21ba_4
XANTENNA__08611__B1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A2 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ net496 net648 _06640_ net417 net1926 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11761__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\] vssd1
+ vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\] vssd1
+ vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ net656 net707 net266 net825 vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold992 team_03_WB.instance_to_wrap.core.register_file.registers_state\[812\] vssd1
+ vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ _03059_ net2028 net288 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10721__A1 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ clknet_leaf_32_wb_clk_i net1929 _01185_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ clknet_leaf_120_wb_clk_i _02515_ _01116_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11963_ net627 _06740_ net465 net369 net2544 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10485__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ clknet_leaf_86_wb_clk_i _01466_ _00067_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__inv_2
X_14682_ clknet_leaf_52_wb_clk_i _02446_ _01047_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11894_ net621 _06703_ net461 net378 net1977 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__a32o_1
XANTENNA__07350__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13633_ net1313 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
X_10845_ net689 _05596_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13564_ net1333 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
X_10776_ net1246 net1015 vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__and2_2
XFILLER_0_54_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11985__A0 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14484__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12515_ net1300 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XANTENNA__07653__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13495_ net1334 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ net1384 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07405__A1 net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15165_ net1546 vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_2
X_12377_ net1353 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
X_14116_ clknet_leaf_19_wb_clk_i _01880_ _00481_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\]
+ sky130_fd_sc_hd__dfrtp_1
X_11328_ _06631_ net2508 net411 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ net1477 vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11259_ net710 _06468_ net822 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__and3_1
X_14047_ clknet_leaf_114_wb_clk_i _01811_ _00412_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[401\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06916__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__B2 _06346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13156__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14949_ clknet_leaf_63_wb_clk_i _02701_ _01314_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08470_ net1055 _04409_ _04410_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07421_ net1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[852\]
+ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07892__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07352_ net1151 _03293_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11976__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__A2 _04775_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07644__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07283_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09022_ net854 _04962_ _04963_ _04961_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__o31a_1
XFILLER_0_2_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold200 _02589_ vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold211 team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\] vssd1
+ vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 team_03_WB.instance_to_wrap.CPU_DAT_I\[22\] vssd1 vssd1 vccd1 vccd1 net1806
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[298\] vssd1
+ vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\] vssd1
+ vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 team_03_WB.instance_to_wrap.core.register_file.registers_state\[7\] vssd1
+ vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold266 team_03_WB.instance_to_wrap.ADR_I\[18\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06988__C_N _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 net184 vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09149__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold288 _02575_ vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 net180 vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ net317 _05863_ _05864_ _05429_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__or4b_1
Xfanout702 _06559_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout713 net715 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1111_A net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1209_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
Xfanout746 net750 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 net759 vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
X_09855_ _05795_ _05796_ _05081_ _05794_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a211o_1
XANTENNA__10703__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A _03024_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 net770 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10703__B2 team_03_WB.instance_to_wrap.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout779 net785 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__buf_2
XANTENNA__11900__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06887__B net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _04744_ _04747_ net865 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o21ai_1
X_09786_ net327 _05384_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a21o_1
X_06998_ _02792_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02939_ vssd1
+ vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ net847 _04663_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_119_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08668_ _04608_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11017__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07332__B1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07619_ net804 _03549_ _03550_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__or3_1
XANTENNA__07883__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _04539_ _04540_ net854 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10630_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] team_03_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ net839 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11967__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07096__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ net2072 net537 net598 _05871_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07635__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07230__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ net1303 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
X_13280_ net1396 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
X_10492_ net2058 net1025 net905 team_03_WB.instance_to_wrap.ADR_I\[14\] vssd1 vssd1
+ vccd1 vccd1 _02617_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ net1695 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11195__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ net1648 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11734__A3 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11113_ net829 _06541_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__and2_2
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _06791_ net462 net447 net2199 vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ net636 _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__nor2_1
X_15069__1450 vssd1 vssd1 vccd1 vccd1 _15069__1450/HI net1450 sky130_fd_sc_hd__conb_1
XANTENNA__07797__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07571__B1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ clknet_leaf_38_wb_clk_i _02567_ _01168_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.BUSY_O
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13724__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12995_ net1296 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11923__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14734_ clknet_leaf_122_wb_clk_i _02498_ _01099_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_11946_ net634 _06723_ net472 net372 net2020 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07323__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09863__A2 _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14665_ clknet_leaf_60_wb_clk_i _02429_ _01030_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ net617 _06686_ net456 net377 net1912 vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11224__A _06456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ net1316 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09076__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10828_ net691 _05499_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__or2_1
XANTENNA__09615__A2 _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14596_ clknet_leaf_17_wb_clk_i _02360_ _00961_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11958__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13547_ net1325 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
XANTENNA__07140__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ _02774_ _06294_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand2_1
XANTENNA__07848__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10630__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__A _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11973__A3 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13478_ net1397 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15217_ net911 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_1
X_12429_ net1290 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11725__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net1529 vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
XFILLER_0_77_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10933__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\]
+ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__or2_1
X_15079_ net1460 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_10_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06988__A team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net873 vssd1 vssd1 vccd1
+ vccd1 _02863_ sky130_fd_sc_hd__and2_4
XANTENNA__09000__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A3 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ _05371_ _05569_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__a21bo_1
X_06852_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[44\] vssd1
+ vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_109_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11118__B _06557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ net577 _05371_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08522_ net937 _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07314__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08511__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[988\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1020\] net1208
+ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10449__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11134__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07404_ net1121 _03342_ _03343_ _03345_ net1131 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a311o_1
XFILLER_0_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ net551 _04296_ _04325_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11949__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07617__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ net721 _03260_ _03269_ _03276_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_50_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10973__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1061_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1159_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07266_ net609 _03205_ _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__o21ai_2
XANTENNA__11964__A3 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\]
+ net954 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07197_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08162__B net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1326_A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__C1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08042__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout786_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 net514 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06898__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07493__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout521 net524 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_8
XANTENNA__09274__A _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
X_09907_ _05541_ _05842_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor2_1
XANTENNA__13747__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout543 _04815_ vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_2
Xfanout554 _03105_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout953_A net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 _03025_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10688__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
X_09838_ net580 _05670_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout587 _06400_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__buf_2
XFILLER_0_57_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07553__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09769_ _04775_ _05106_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net2427 _06519_ net333 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__mux2_1
XANTENNA__13897__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ net1303 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07305__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10867__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ net593 _06505_ net469 _06808_ net1795 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a32o_1
XFILLER_0_132_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14450_ clknet_leaf_101_wb_clk_i _02214_ _00815_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ net2607 _06625_ net352 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__mux2_1
XANTENNA__09058__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13401_ net1309 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XANTENNA__07608__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ net1671 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] net835 vssd1 vssd1 vccd1
+ vccd1 _02515_ sky130_fd_sc_hd__mux2_1
X_11593_ net271 net2407 net452 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__mux2_1
X_14381_ clknet_leaf_105_wb_clk_i _02145_ _00746_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10883__A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ team_03_WB.instance_to_wrap.WRITE_I team_03_WB.instance_to_wrap.READ_I vssd1
+ vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input82_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13332_ net1321 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XANTENNA__11955__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08353__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10475_ net2054 net1026 net902 team_03_WB.instance_to_wrap.ADR_I\[31\] vssd1 vssd1
+ vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
X_13263_ net1390 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15002_ clknet_leaf_23_wb_clk_i net50 _01367_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14522__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ net1606 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13194_ net1256 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10107__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12145_ net1718 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11918__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12076_ _06782_ net464 net444 net1801 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ net704 net271 net823 vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__and3_1
XANTENNA__11340__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__A _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11653__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12978_ net1420 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07432__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ clknet_leaf_120_wb_clk_i _02481_ _01082_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11929_ _06505_ net2766 net375 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09049__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14648_ clknet_leaf_10_wb_clk_i _02412_ _01013_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14579_ clknet_leaf_115_wb_clk_i _02343_ _00944_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[933\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ net722 _03058_ _03043_ net612 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11946__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07051_ net611 _02989_ _02991_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08024__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07953_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\] net788
+ _03892_ net1145 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__o211a_1
XANTENNA__08202__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ net1132 net898 vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nor2_8
XANTENNA__11129__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\]
+ net899 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07535__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09623_ _05482_ _05494_ net572 vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__mux2_1
X_06835_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 _02778_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout367_A net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ net325 _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06884__C team_03_WB.instance_to_wrap.core.decoder.inst\[27\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08505_ net544 net440 net429 _04444_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__or4_1
X_09485_ net325 _05419_ _05422_ net584 _05426_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__a221o_1
XANTENNA__11634__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10842__A0 _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1276_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_77_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08367_ _04303_ _04308_ net867 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout701_A _06559_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07318_ net812 _03258_ _03259_ _03251_ _03254_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a32o_1
XANTENNA__14545__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09269__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[184\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\] net984 net925
+ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07249_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[168\]
+ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _06098_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__nor2_1
XANTENNA__09212__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09763__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] net672 vssd1 vssd1 vccd1
+ vccd1 _06033_ sky130_fd_sc_hd__nand2_1
XANTENNA__10642__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1305 net1317 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__buf_2
XFILLER_0_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1316 net1317 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__clkbuf_4
Xfanout1327 net1328 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1338 net1339 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__buf_4
Xfanout340 _06809_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__buf_4
Xfanout1349 net1359 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__clkbuf_2
Xfanout351 net352 vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__buf_4
Xfanout362 _06818_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_4
X_13950_ clknet_leaf_58_wb_clk_i _01714_ _00315_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[304\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_6
Xfanout384 _06812_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07526__B1 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_8
X_12901_ net1277 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
X_13881_ clknet_leaf_93_wb_clk_i _01645_ _00246_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07541__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ net1408 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09818__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12763_ net1348 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11625__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14502_ clknet_leaf_78_wb_clk_i _02266_ _00867_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[856\]
+ sky130_fd_sc_hd__dfrtp_1
X_11714_ net2257 _06418_ net341 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__mux2_1
XANTENNA__10833__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ net1345 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14433_ clknet_leaf_1_wb_clk_i _02197_ _00798_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10817__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11645_ net2430 _06611_ net348 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14364_ clknet_leaf_125_wb_clk_i _02128_ _00729_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[718\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08083__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_1
X_11576_ net281 net2704 net454 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
Xinput37 gpio_in[12] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10597__C1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput48 gpio_in[23] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput59 gpio_in[34] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XANTENNA__10061__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13912__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ net1289 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
X_10527_ net139 net1023 net1019 net1873 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ clknet_leaf_87_wb_clk_i _02059_ _00660_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[649\]
+ sky130_fd_sc_hd__dfrtp_1
X_10458_ _06272_ _06271_ net284 vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__mux2_1
XANTENNA__09907__A _05541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13246_ net1414 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11648__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10389_ _05994_ _05995_ _06085_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__and3_1
XANTENNA__11875__C net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13177_ net1352 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XANTENNA__07765__B1 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08962__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net1697 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09506__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12059_ _06625_ net2699 net362 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08714__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09809__A2 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11616__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ net588 _05210_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08493__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09690__B1 _05631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08221_ _04157_ _04162_ net871 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08152_ net850 _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08245__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07048__A2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07103_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\]
+ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__and2_1
XFILLER_0_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11131__B net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07453__C1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__or3_1
XANTENNA__10052__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07034_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\]
+ net895 vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06940__S net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07205__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1024_A _06283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09028__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08985_ _04925_ _04926_ net851 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A3 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\] net1146
+ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07508__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14098__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07867_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[347\]
+ net780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\] net1127
+ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout749_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13074__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ _05546_ _05547_ net578 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07798_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__or3_1
XANTENNA__07072__A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ net591 _05456_ _05457_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__o31a_1
XFILLER_0_116_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout916_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10815__B1 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ net561 _05101_ _05103_ _05409_ net571 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__o311a_1
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07800__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ net851 _04359_ _04360_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or3_1
XFILLER_0_136_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10637__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _03352_ _04475_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09659__S1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11430_ net506 _06537_ _06756_ net403 net1994 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a32o_1
XANTENNA__08236__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ net1241 net832 _06477_ net666 vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__and4_1
XFILLER_0_116_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ team_03_WB.instance_to_wrap.core.pc.current_pc\[31\] _06153_ vssd1 vssd1
+ vccd1 vccd1 _06154_ sky130_fd_sc_hd__xnor2_1
X_13100_ net1298 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
XANTENNA__11791__A1 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14080_ clknet_leaf_130_wb_clk_i _01844_ _00445_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\]
+ sky130_fd_sc_hd__dfrtp_1
X_11292_ net511 net637 _06713_ net415 net2244 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ net1403 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
X_10243_ _05999_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__or2_1
XANTENNA__11543__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08944__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] net821 _06015_ vssd1
+ vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A gpio_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 net1105 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
Xfanout1113 net1114 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1124 net1125 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_4
Xfanout1135 net1136 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14982_ clknet_leaf_124_wb_clk_i net61 _01347_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12099__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1157 net1160 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_4
Xfanout1168 net1198 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06970__A1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06970__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13933_ clknet_leaf_110_wb_clk_i _01697_ _00298_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10401__A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13864_ clknet_leaf_26_wb_clk_i _01628_ _00229_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08078__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ net1380 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13795_ clknet_leaf_21_wb_clk_i _01559_ _00160_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11931__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ net1249 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12677_ net1275 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06858__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08227__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416_ clknet_leaf_80_wb_clk_i _02180_ _00781_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\]
+ sky130_fd_sc_hd__dfrtp_1
X_11628_ _06702_ net387 net356 net2529 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11231__A0 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ clknet_leaf_45_wb_clk_i _02111_ _00712_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11559_ net655 _06669_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__nor2_1
XANTENNA__10585__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold607 team_03_WB.instance_to_wrap.core.register_file.registers_state\[642\] vssd1
+ vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\] vssd1
+ vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold629 team_03_WB.instance_to_wrap.core.register_file.registers_state\[825\] vssd1
+ vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ clknet_leaf_74_wb_clk_i _02042_ _00643_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13229_ net1319 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__B_N _03489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08770_ net441 net433 _04711_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__or3_2
XANTENNA__08687__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09372__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ net1109 _03661_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor3_1
XANTENNA__11298__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11837__A2 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08163__B1 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07652_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[846\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\] net1145
+ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11126__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07583_ net1141 _03514_ _03524_ net722 vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_88_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09322_ _04711_ _05255_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__xor2_1
XANTENNA__08466__A1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07958__A1_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06935__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10965__B _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11470__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07674__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _03604_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ net867 _04137_ _04140_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ net579 net572 _05124_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__and3_1
XANTENNA__12014__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11222__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ _03641_ _03823_ _04031_ _04071_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__B1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__A1 net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07017_ net1125 _02956_ _02957_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1406_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07067__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[713\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[745\] net941
+ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07919_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\] net782
+ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11828__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ net851 _04839_ _04840_ _04838_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10930_ net690 _06515_ _06516_ _06514_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__a31o_4
Xclkbuf_leaf_92_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10500__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14883__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10861_ net1240 _06388_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__o21a_2
XFILLER_0_6_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09103__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net1370 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XANTENNA__08457__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13580_ net1310 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10792_ net684 net315 vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XANTENNA__07530__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ net1264 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10803__A3 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ net1338 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14201_ clknet_leaf_83_wb_clk_i _01965_ _00566_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11413_ _06478_ _06751_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15181_ net1562 vssd1 vssd1 vccd1 vccd1 la_data_out[117] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12393_ net1252 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10567__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07968__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ clknet_leaf_90_wb_clk_i _01896_ _00497_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11344_ net503 net624 _06724_ net406 net2377 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a32o_1
XFILLER_0_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09709__A1 _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14063_ clknet_leaf_102_wb_clk_i _01827_ _00428_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ net712 _06504_ net824 vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__and3_1
X_13014_ net1345 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09185__A2 _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ _06006_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or2_1
XANTENNA__07196__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _03943_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 team_03_WB.instance_to_wrap.core.register_file.registers_state\[952\] vssd1
+ vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14965_ clknet_leaf_55_wb_clk_i _02717_ _01330_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ net591 _05456_ _05457_ _05478_ _05499_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__o311a_1
XANTENNA__11819__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13916_ clknet_leaf_129_wb_clk_i _01680_ _00281_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07043__S1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14896_ clknet_leaf_45_wb_clk_i _02659_ _01261_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09893__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ clknet_leaf_72_wb_clk_i _01611_ _00212_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11661__S net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08448__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13778_ clknet_leaf_101_wb_clk_i _01542_ _00143_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12729_ net1356 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07120__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15191__1572 vssd1 vssd1 vccd1 vccd1 _15191__1572/HI net1572 sky130_fd_sc_hd__conb_1
XFILLER_0_127_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11204__A0 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10558__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold404 _02600_ vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold415 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\] vssd1
+ vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15208__1576 vssd1 vssd1 vccd1 vccd1 _15208__1576/HI net1576 sky130_fd_sc_hd__conb_1
Xhold426 team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\] vssd1
+ vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\] vssd1
+ vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 team_03_WB.instance_to_wrap.CPU_DAT_I\[8\] vssd1 vssd1 vccd1 vccd1 net2032
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09940_ _05874_ net2136 net293 vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__mux2_1
XANTENNA__07974__A3 net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold459 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\] vssd1
+ vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
X_09871_ _05198_ _05634_ net591 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a21o_1
Xfanout917 net919 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_4
Xfanout928 _04088_ vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_2
XANTENNA__07187__A1 net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout939 net945 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
X_08822_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\] net1000 net1204
+ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__o221a_1
XANTENNA__08923__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10740__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\] vssd1
+ vssd1 vccd1 vccd1 net2688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\] vssd1
+ vssd1 vccd1 vccd1 net2699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06934__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1126 team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\] vssd1
+ vssd1 vccd1 vccd1 net2710 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07615__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\] vssd1
+ vssd1 vccd1 vccd1 net2721 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\] net976
+ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__or2_1
Xhold1148 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\] vssd1
+ vssd1 vccd1 vccd1 net2732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13780__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1159 team_03_WB.instance_to_wrap.core.register_file.registers_state\[152\] vssd1
+ vssd1 vccd1 vccd1 net2743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07704_ net741 _03642_ _03643_ _03644_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__o32a_1
XFILLER_0_75_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08684_ _04622_ _04623_ _04624_ _04625_ net860 net922 vssd1 vssd1 vccd1 vccd1 _04626_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09884__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07635_ net801 _03572_ _03575_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__a22o_1
XANTENNA__11691__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07895__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1189_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ net1191 team_03_WB.instance_to_wrap.core.register_file.registers_state\[728\]
+ net777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\] net745
+ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ net607 _05144_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07647__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07497_ _03437_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout1356_A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09976__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07662__A2 _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14286__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09167_ net443 net435 _04953_ net554 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08118_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[986\]
+ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ net863 _05039_ _05034_ net846 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout983_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08049_ net1178 team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\]
+ net874 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\] vssd1
+ vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold971 team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\] vssd1
+ vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold982 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\] vssd1
+ vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11060_ net2660 net426 _06607_ net511 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
Xhold993 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\] vssd1
+ vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10011_ _03023_ net1813 net291 vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10650__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12431__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11047__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ clknet_leaf_40_wb_clk_i _02514_ _01115_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11962_ net632 _06739_ net470 net371 net2242 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09875__B1 _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ clknet_leaf_107_wb_clk_i _01465_ _00066_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10913_ net690 _06501_ _06502_ _06500_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a31o_4
X_14681_ clknet_leaf_52_wb_clk_i _02445_ _01046_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11682__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ net627 _06702_ net465 net378 net2309 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ net1330 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
X_10844_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[21\] net309 net689 vssd1
+ vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__a21o_1
XANTENNA__11434__A0 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13563_ net1310 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10775_ _02930_ _06384_ _06383_ _02942_ _02934_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ net1346 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08790__S net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13494_ net1334 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12445_ net1382 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XANTENNA__11737__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12606__A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14779__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08063__C1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08602__A1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15164_ net1545 vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08091__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ net1362 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14115_ clknet_leaf_24_wb_clk_i _01879_ _00480_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\]
+ sky130_fd_sc_hd__dfrtp_1
X_11327_ net264 net2709 net412 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__mux2_1
X_15095_ net1476 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
X_14046_ clknet_leaf_57_wb_clk_i _01810_ _00411_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09915__A _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ net495 net619 _06696_ net413 net2352 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a32o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11656__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ _06043_ _06050_ _06042_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10173__A0 _04954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12341__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net510 net654 _06675_ net419 net1828 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14948_ clknet_leaf_30_wb_clk_i _02700_ _01313_ vssd1 vssd1 vccd1 vccd1 team_03_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11268__A3 _06701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10476__B2 team_03_WB.instance_to_wrap.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07877__C1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14879_ clknet_leaf_51_wb_clk_i _02642_ _01244_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07341__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07420_ _03355_ _03356_ _03361_ net1151 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07629__C1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\]
+ net757 net1115 vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__mux4_1
XFILLER_0_50_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09633__A3 _05570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A2 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07282_ net819 _03222_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10087__A_N _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09021_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[208\]
+ net981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\] net944
+ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11420__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08054__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 net215 vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 net195 vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 _02593_ vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 net237 vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold245 team_03_WB.instance_to_wrap.CPU_DAT_I\[1\] vssd1 vssd1 vccd1 vccd1 net1829
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold256 team_03_WB.instance_to_wrap.core.register_file.registers_state\[418\] vssd1
+ vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _02621_ vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 team_03_WB.instance_to_wrap.CPU_DAT_I\[11\] vssd1 vssd1 vccd1 vccd1 net1862
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10951__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09923_ _05863_ _05864_ net314 _05429_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__and4bb_2
Xhold289 team_03_WB.instance_to_wrap.CPU_DAT_I\[12\] vssd1 vssd1 vccd1 vccd1 net1873
+ sky130_fd_sc_hd__dlygate4sd3_1
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout714 net715 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout397_A net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net728 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
Xfanout736 _02853_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_4
Xfanout747 net750 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__clkbuf_4
X_09854_ net569 _05792_ _05793_ net580 vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__o31a_1
Xfanout758 net759 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1104_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09036__S net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ net860 _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__and3_1
XANTENNA__07345__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09785_ _03459_ _04619_ _04820_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08109__B1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ _02927_ _02929_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08736_ net1077 _04670_ _04677_ net843 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07868__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\] net1074
+ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a221o_1
XANTENNA__07332__A1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _03558_ _03559_ net810 vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a21o_1
X_15118__1499 vssd1 vssd1 vccd1 vccd1 _15118__1499/HI net1499 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07883__A2 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\] net920
+ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11416__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07549_ _03459_ _03489_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10560_ net2197 net534 net595 _05870_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XANTENNA__14921__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ net605 _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nor2_1
XANTENNA__10645__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ net1967 net1025 net905 team_03_WB.instance_to_wrap.ADR_I\[15\] vssd1 vssd1
+ vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11719__A1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12230_ net1742 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08045__C1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07399__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11195__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ net1592 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07954__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11112_ net264 net2619 net422 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__mux2_1
X_12092_ _06790_ net461 net447 net1993 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a22o_1
Xhold790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\] vssd1
+ vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11043_ net712 _06517_ net702 vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08899__A1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15190__1571 vssd1 vssd1 vccd1 vccd1 _15190__1571/HI net1571 sky130_fd_sc_hd__conb_1
XANTENNA__07571__A1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ clknet_leaf_56_wb_clk_i _02566_ _01167_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ net1366 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ clknet_leaf_15_wb_clk_i _02497_ _01098_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14451__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ net617 _06722_ net456 net369 net2826 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14664_ clknet_leaf_33_wb_clk_i _02428_ _01029_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1018\]
+ sky130_fd_sc_hd__dfstp_1
X_11876_ net631 _06685_ net471 net380 net2064 vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11407__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13615_ net1421 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
X_10827_ net277 net2268 net523 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XANTENNA__09076__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14595_ clknet_leaf_25_wb_clk_i _02359_ _00960_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[949\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13546_ net1325 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
XANTENNA__12080__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ net1932 net532 net527 _06372_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a22o_1
XANTENNA__08823__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13477_ net1397 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
XANTENNA__09629__B _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ _05563_ _06312_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or2_1
XANTENNA__12336__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15216_ net910 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_1
X_12428_ net1300 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ net1528 vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
XFILLER_0_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12359_ net1390 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10933__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15078_ net1459 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_43_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14029_ clknet_leaf_104_wb_clk_i _01793_ _00394_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\]
+ sky130_fd_sc_hd__dfrtp_1
X_06920_ _02858_ _02861_ net814 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09000__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__B2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11894__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _02794_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09570_ net325 _05378_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08521_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[191\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\] net971 net920
+ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08511__B1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07403_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1023\]
+ net893 _03344_ net1147 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o311a_1
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11134__B net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08383_ net437 net429 _04323_ net544 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07078__B1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ net812 _03275_ net717 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06943__S net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10621__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07265_ net612 _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08443__B _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A _02791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\] net914
+ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07196_ net1200 net1012 _03107_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__a21o_1
XANTENNA__08578__B1 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11177__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1221_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1319_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07250__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 net505 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout779_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout511 net514 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
X_09906_ _05596_ _05833_ _05847_ _05500_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or4b_1
Xfanout522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_6
Xfanout533 _06309_ vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout544 net546 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__buf_2
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10688__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 _03025_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07075__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ net569 _05721_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__nand2_1
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14474__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 _06299_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_2
XANTENNA_fanout946_A net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09768_ _05092_ _05120_ net579 vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08719_ net1214 _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__and3_1
XANTENNA__11637__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07305__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _04816_ _05639_ net664 vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11730_ net1980 _06499_ net341 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07856__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09058__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ net2202 _06624_ net352 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__mux2_1
XANTENNA__07241__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ net1308 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ net2421 net2878 net835 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__mux2_1
XANTENNA__07069__B1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380_ clknet_leaf_6_wb_clk_i _02144_ _00745_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[734\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _06487_ net2500 net455 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13331_ net1330 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10543_ net1792 net1024 net905 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input75_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13262_ net1282 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XANTENNA__08018__C1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ net1 net1024 vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15001_ clknet_leaf_124_wb_clk_i net49 _01366_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ net1605 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13193_ net1251 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12144_ net1658 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12075_ _06781_ net460 net444 net2142 vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11026_ net2776 net426 _06587_ net518 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a22o_1
XANTENNA__09533__A2 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11876__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07416__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08741__B1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07544__B2 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__B _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11891__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07713__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11628__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ net1305 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
XANTENNA__11235__A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ clknet_leaf_116_wb_clk_i _02480_ _01081_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_11928_ _06626_ net2847 net373 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09049__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14647_ clknet_leaf_76_wb_clk_i _02411_ _01012_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1001\]
+ sky130_fd_sc_hd__dfstp_1
X_11859_ net300 net2822 net383 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12053__A0 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08257__C1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ clknet_leaf_100_wb_clk_i _02342_ _00943_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_138_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08544__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10603__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13529_ net1327 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07050_ net611 _02989_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a21o_1
XANTENNA__07480__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_109_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_122_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_50_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10906__A2 _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_2_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
X_15117__1498 vssd1 vssd1 vccd1 vccd1 _15117__1498/HI net1498 sky130_fd_sc_hd__conb_1
X_07952_ net1140 _03884_ _03885_ _03893_ net1157 vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o311a_1
XANTENNA__12005__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ net1014 net1012 net1015 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11867__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11129__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ net1192 net880 team_03_WB.instance_to_wrap.core.register_file.registers_state\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a21o_1
XANTENNA__07535__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ _05331_ _05335_ _05337_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or3_1
X_06834_ team_03_WB.instance_to_wrap.READ_I vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06938__S net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08719__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11882__A3 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _05493_ _05494_ net566 vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__mux2_1
XANTENNA__11619__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08504_ _04080_ _04444_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nor2_1
XANTENNA__08496__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _05425_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[922\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13360__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1269_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08366_ net1210 _04306_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07317_ net802 _03247_ _03248_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08297_ net941 _04238_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09984__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07471__B1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07248_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[8\] net774
+ net747 _03189_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout896_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09212__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ net1151 _03119_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10190_ _06030_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__nand2_1
XANTENNA__07774__A1 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1306 net1307 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__buf_4
Xfanout1317 net1433 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__clkbuf_4
Xfanout1328 net1335 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_6
Xfanout1339 net1359 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__buf_2
Xfanout341 net343 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_6
XANTENNA__11858__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout352 _06805_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_4
Xfanout363 net364 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_8
Xfanout374 _06814_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_4
XANTENNA__07526__A1 net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 net387 vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_4
X_12900_ net1311 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
Xfanout396 _06778_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_8
X_13880_ clknet_leaf_8_wb_clk_i _01644_ _00245_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10530__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12831_ net1378 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12762_ net1370 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ clknet_leaf_108_wb_clk_i _02265_ _00866_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ net1890 _06413_ net341 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12693_ net1268 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14432_ clknet_leaf_132_wb_clk_i _02196_ _00797_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12035__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11644_ net2442 _06609_ net351 vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14363_ clknet_leaf_28_wb_clk_i _02127_ _00728_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ _06390_ _06394_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__nand2_4
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 gpio_in[13] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ net1289 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10526_ net140 net1023 net1019 net1928 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
Xinput49 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ clknet_leaf_83_wb_clk_i _02058_ _00659_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11929__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13245_ net1381 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
X_10457_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] _06134_ vssd1 vssd1 vccd1
+ vccd1 _06272_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09907__B _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08411__C1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net1369 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
X_10388_ _05994_ _05995_ _06085_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07765__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08962__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ net1657 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06973__C1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ _06624_ net2527 net362 vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__mux2_1
XANTENNA__07517__A1 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08714__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11664__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net624 _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__nor2_1
XANTENNA__10521__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08478__C1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10824__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09690__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ net1212 _04160_ _04161_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__o21a_1
XANTENNA__13180__A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12026__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13737__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08151_ net1220 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\]
+ net949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\] net929
+ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07102_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[417\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[385\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[289\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[257\]
+ net776 net1123 vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux4_1
XANTENNA__07453__B1 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10052__A2 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08082_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\] net789
+ net1011 _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10028__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07033_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\] net776
+ net746 _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08402__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07756__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ net1223 team_03_WB.instance_to_wrap.core.register_file.registers_state\[138\]
+ net957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[170\] net931
+ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout1017_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07935_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\] vssd1
+ vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__o22a_1
XANTENNA__09053__S0 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07866_ net1158 _03807_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__nor2_1
XANTENNA__10512__B1 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08181__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _05459_ _05466_ net574 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__mux2_1
XANTENNA__08181__B2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07353__A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07797_ _03731_ _03732_ _03737_ _03738_ net1111 net1131 vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout644_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1386_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__inv_2
XANTENNA__10815__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ net561 _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__nand2_1
XANTENNA__09681__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13090__A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08418_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[218\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\] net933
+ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o221a_1
XANTENNA__12017__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09398_ _05170_ _05174_ _05338_ _05172_ _05167_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_65_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net1056 _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__or3_1
XANTENNA__10579__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11240__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ net494 net616 _06732_ net405 net2209 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08912__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06152_ vssd1 vssd1
+ vccd1 vccd1 _06153_ sky130_fd_sc_hd__nand2_1
XANTENNA__10653__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ net715 _06541_ net824 vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__and3_1
XANTENNA__08619__S0 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13030_ net1423 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
X_10242_ _06080_ _06081_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08944__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _04954_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] net673 vssd1
+ vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__mux2_1
Xfanout1103 net1105 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1114 _02786_ vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06955__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1125 net1129 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_2
Xfanout1136 team_03_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_A gpio_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 team_03_WB.instance_to_wrap.core.decoder.inst\[22\] vssd1 vssd1 vccd1
+ vccd1 net1147 sky130_fd_sc_hd__clkbuf_8
Xfanout1158 net1159 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_8
X_14981_ clknet_leaf_124_wb_clk_i net34 _01346_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1169 net1170 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_2
XANTENNA__13265__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13932_ clknet_leaf_9_wb_clk_i _01696_ _00297_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08172__A1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ clknet_leaf_69_wb_clk_i _01627_ _00228_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[217\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12814_ net1336 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
XANTENNA__14192__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ clknet_leaf_131_wb_clk_i _01558_ _00159_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[148\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__A1_N team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12745_ net1247 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116__1497 vssd1 vssd1 vccd1 vccd1 _15116__1497/HI net1497 sky130_fd_sc_hd__conb_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12008__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ net1311 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
X_14415_ clknet_leaf_99_wb_clk_i _02179_ _00780_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[769\]
+ sky130_fd_sc_hd__dfrtp_1
X_11627_ _06701_ net390 net354 net2513 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12023__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10034__A2 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09918__A _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07435__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14346_ clknet_leaf_10_wb_clk_i _02110_ _00711_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08632__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ net2279 net489 _06793_ net517 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11659__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\] vssd1
+ vssd1 vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10509_ net159 net1023 net1019 net2037 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
Xhold619 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\] vssd1
+ vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
X_14277_ clknet_leaf_108_wb_clk_i _02041_ _00642_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11489_ _06609_ net2791 net396 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13228_ net1299 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08935__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ net1401 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07720_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\] net726
+ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__o221a_1
XANTENNA__11298__A1 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11837__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07173__A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ net751 _03590_ _03592_ net1107 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07910__A1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15049__1581 vssd1 vssd1 vccd1 vccd1 net1581 _15049__1581/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ net1159 _03519_ _03521_ _03523_ net1132 vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10030__C net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09321_ _05260_ _05261_ _05259_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__a21o_1
XANTENNA__10738__S net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11470__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _03728_ _05147_ net606 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07674__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08203_ _04141_ _04142_ _04143_ _04144_ net855 net930 vssd1 vssd1 vccd1 vccd1 _04145_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09183_ net572 _05124_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08134_ _03459_ _03489_ _03280_ _03314_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10981__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ net812 _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09179__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[835\]
+ net1148 vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a21o_1
XANTENNA__07729__A1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11525__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1301_A net1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10733__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[617\] net925
+ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07918_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\]
+ net880 _02872_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\] net917
+ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07849_ net1192 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\]
+ net883 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__and3_1
XANTENNA__07901__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10860_ net1039 net1245 net1246 _02808_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__or4_4
XFILLER_0_116_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__B1 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ net568 _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__nand2_1
XANTENNA__09654__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _02829_ net688 _06399_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12530_ net1398 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11333__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ net1268 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14200_ clknet_leaf_10_wb_clk_i _01964_ _00565_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[554\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ _06473_ net2712 net401 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15180_ net1561 vssd1 vssd1 vccd1 vccd1 la_data_out[116] sky130_fd_sc_hd__buf_2
XANTENNA__09738__A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12392_ net1285 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
XANTENNA__08614__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07968__A1 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07512__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ clknet_leaf_111_wb_clk_i _01895_ _00496_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[485\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11343_ net1242 net832 net278 net666 vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10972__B1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__A2 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ clknet_leaf_72_wb_clk_i _01826_ _00427_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\]
+ sky130_fd_sc_hd__dfrtp_1
X_11274_ net501 net622 _06704_ net413 net2370 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ net1262 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
X_10225_ _06008_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08393__A1 net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _04984_ net674 _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold5 team_03_WB.instance_to_wrap.core.register_file.registers_state\[940\] vssd1
+ vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
X_14964_ clknet_leaf_56_wb_clk_i _02716_ _01329_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10087_ _05686_ _05697_ _05706_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13915_ clknet_leaf_35_wb_clk_i _01679_ _00280_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14895_ clknet_leaf_37_wb_clk_i _02658_ _01260_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09920__B _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13846_ clknet_leaf_82_wb_clk_i _01610_ _00211_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[200\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07721__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09412__S _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13777_ clknet_leaf_95_wb_clk_i _01541_ _00142_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07105__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ net280 net648 net703 net822 vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__and4_1
XANTENNA__08536__B _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11243__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07656__B1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__D_N _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08853__C1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12728_ net1368 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07120__A2 _03058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12659_ net1266 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09648__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07959__A1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold405 net116 vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14329_ clknet_leaf_112_wb_clk_i _02093_ _00694_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold416 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\] vssd1
+ vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold427 team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\] vssd1
+ vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold438 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\] vssd1
+ vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 net207 vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08908__B1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__inv_2
XANTENNA__09176__A3 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout907 _05907_ vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09030__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout929 net930 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_4
X_08821_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\] net1000
+ _04762_ net1072 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__o211a_1
Xhold1105 team_03_WB.instance_to_wrap.core.register_file.registers_state\[585\] vssd1
+ vssd1 vccd1 vccd1 net2689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1116 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\] vssd1
+ vssd1 vccd1 vccd1 net2700 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\] vssd1
+ vssd1 vccd1 vccd1 net2711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08752_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[643\] net976 vssd1
+ vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__a22o_1
Xhold1138 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\] vssd1
+ vssd1 vccd1 vccd1 net2722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 team_03_WB.instance_to_wrap.core.register_file.registers_state\[664\] vssd1
+ vssd1 vccd1 vccd1 net2733 sky130_fd_sc_hd__dlygate4sd3_1
X_07703_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\]
+ net891 net1120 vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08683_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__mux2_1
XANTENNA__11852__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07344__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07634_ net742 _03574_ net806 vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07631__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10468__S net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ net1188 team_03_WB.instance_to_wrap.core.register_file.registers_state\[600\]
+ net777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[632\] net732
+ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o221a_1
XFILLER_0_7_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1084_A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09100__A3 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15159__1540 vssd1 vssd1 vccd1 vccd1 _15159__1540/HI net1540 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07496_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\] net733
+ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09235_ _04235_ _05175_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10992__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1251_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A _02938_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1349_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ net443 net435 _04893_ net547 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08117_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\]
+ net891 _04058_ net1119 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__o311a_1
XANTENNA__11746__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09097_ _05035_ _05036_ _05038_ _05037_ net933 net858 vssd1 vssd1 vccd1 vccd1 _05039_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08611__A2 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08048_ _03945_ _03946_ _03986_ _03987_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__o22a_1
Xhold950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\] vssd1
+ vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\] vssd1
+ vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout976_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold972 team_03_WB.instance_to_wrap.core.register_file.registers_state\[919\] vssd1
+ vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold983 net154 vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09167__A3 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[778\] vssd1
+ vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ net590 net1755 net289 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15115__1496 vssd1 vssd1 vccd1 vccd1 _15115__1496/HI net1496 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _05884_ net1785 net290 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07583__C1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08127__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11961_ net622 _06738_ net462 net370 net2366 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09875__B2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ net315 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__or4b_1
X_13700_ clknet_leaf_15_wb_clk_i _01464_ _00065_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_14680_ clknet_leaf_52_wb_clk_i _02444_ _01045_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11892_ net641 _06701_ net481 net379 net2201 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13631_ net1400 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10843_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[21\] net307 vssd1
+ vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11063__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ net1310 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
X_10774_ _02831_ _02838_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12513_ net1287 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13493_ net1334 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12444_ net1355 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15163_ net1544 vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12375_ net1414 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14380__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14114_ clknet_leaf_130_wb_clk_i _01878_ _00479_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[468\]
+ sky130_fd_sc_hd__dfrtp_1
X_11326_ _06630_ net2636 net412 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15094_ net1475 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13948__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ clknet_leaf_60_wb_clk_i _01809_ _00410_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\]
+ sky130_fd_sc_hd__dfrtp_1
X_11257_ _06453_ net710 net822 vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__and3_1
XANTENNA__09915__B _05676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08366__A1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10208_ _06047_ _06048_ _06046_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ net1040 net833 _06536_ net667 vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__and4_2
XFILLER_0_101_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11370__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _03390_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09931__A _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14947_ clknet_leaf_38_wb_clk_i _00009_ _01312_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11672__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11673__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ clknet_leaf_50_wb_clk_i _02641_ _01243_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07341__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07451__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ clknet_leaf_107_wb_clk_i _01593_ _00194_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07629__B1 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\]
+ net757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08826__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11425__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07281_ net748 _03220_ _03221_ net803 vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\]
+ net981 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\] net928
+ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o221a_1
XANTENNA__14723__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11189__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11420__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08054__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 net227 vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 team_03_WB.instance_to_wrap.CPU_DAT_I\[20\] vssd1 vssd1 vccd1 vccd1 net1797
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\] vssd1
+ vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\] vssd1
+ vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold246 _02572_ vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07329__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold257 team_03_WB.instance_to_wrap.CPU_DAT_I\[23\] vssd1 vssd1 vccd1 vccd1 net1841
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11847__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14873__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold268 team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\] vssd1
+ vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13628__A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold279 _02582_ vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _05517_ _05541_ _05563_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09003__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 _06461_ vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__clkbuf_4
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08357__A1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07626__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout737 net738 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
X_09853_ net567 _05738_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__nand2_1
XANTENNA__08221__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 net750 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07565__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11148__A _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[193\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\] net923
+ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a221o_1
X_09784_ _03459_ _04619_ _05725_ _02945_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__o22a_1
XANTENNA__08109__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06996_ _02925_ _02927_ _02932_ _02934_ _02926_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_77_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08735_ _04674_ _04676_ team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1
+ vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__o21a_1
XANTENNA__10987__A net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__S net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1299_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11664__A1 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[665\]
+ net733 _03547_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\] net937
+ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__S net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__inv_2
XANTENNA__08817__C1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07096__A1 net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07479_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[789\] net789
+ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10926__S net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09218_ _03823_ _05143_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09288__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ net110 net1025 net905 net1897 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ net546 _04296_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10927__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ net1640 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08920__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09749__B1_N net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ _06630_ net2695 net423 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
X_12091_ net620 _06659_ net459 net444 net1779 vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__a32o_1
XANTENNA__10661__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold780 team_03_WB.instance_to_wrap.core.register_file.registers_state\[352\] vssd1
+ vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\] vssd1
+ vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ net2250 net426 _06597_ net516 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07556__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ clknet_leaf_32_wb_clk_i _02565_ _01166_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09848__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07308__C1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ net1268 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XANTENNA__11492__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14732_ clknet_leaf_46_wb_clk_i _02496_ _01097_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11655__A1 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11944_ net629 _06721_ net467 net369 net1888 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a32o_1
XFILLER_0_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14663_ clknet_leaf_63_wb_clk_i _02427_ _01028_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\]
+ sky130_fd_sc_hd__dfstp_1
X_11875_ net1040 net658 net702 net472 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13614_ net1430 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10826_ _06427_ _06429_ net587 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__o21a_2
XANTENNA__14746__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14594_ clknet_leaf_129_wb_clk_i _02358_ _00959_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\]
+ sky130_fd_sc_hd__dfstp_1
X_10757_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] _05769_ net602 vssd1
+ vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__mux2_1
X_13545_ net1281 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13476_ net1397 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ net525 _06327_ _06328_ net530 net2865 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07210__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13770__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15215_ net1579 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
X_12427_ net1253 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08036__B1 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15146_ net1527 vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
X_12358_ net1416 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XANTENNA__11591__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__S net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10933__A3 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ _06619_ net2603 net409 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__mux2_1
X_15077_ net1458 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
X_12289_ net1287 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14028_ clknet_leaf_5_wb_clk_i _01792_ _00393_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06850_ net1244 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__inv_2
XANTENNA__11894__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09839__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08520_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[63\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[31\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
XANTENNA__13183__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07314__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ _04391_ _04392_ net863 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07402_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[991\]
+ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08382_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11134__C net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07333_ net1153 _03273_ _03274_ _03270_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07078__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15114__1495 vssd1 vssd1 vccd1 vccd1 _15114__1495/HI net1495 sky130_fd_sc_hd__conb_1
XFILLER_0_2_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_118_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07264_ team_03_WB.instance_to_wrap.core.decoder.inst\[28\] net821 vssd1 vssd1 vccd1
+ vccd1 _03206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09003_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\] net931
+ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a221o_1
XANTENNA__11150__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ _03108_ _03136_ net610 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__mux2_2
XFILLER_0_103_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout305_A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11582__A0 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11577__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1214_A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout501 net504 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09905_ _05611_ _05623_ _05632_ _05812_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nand4_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 net514 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_4
Xfanout523 net524 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_6
Xfanout534 net538 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14619__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net546 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_1
XANTENNA__11334__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout556 _03064_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_4
XANTENNA__07002__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ net558 _04713_ _05777_ net569 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__a211o_1
XANTENNA__11885__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 net569 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout578 _02993_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_2
XANTENNA__07553__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06979_ net723 _02906_ _02913_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__o22a_4
X_09767_ _05707_ _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout841_A net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__S0 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[420\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[388\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[292\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[260\]
+ net975 net1073 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__mux4_1
X_09698_ _02804_ _03864_ _04820_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07091__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08649_ _04579_ _04590_ net847 vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__mux2_4
XFILLER_0_138_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07710__C1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11660_ net2349 _06623_ net349 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10611_ net1740 net2867 net836 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ net272 net2473 net455 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__mux2_1
XANTENNA__10656__S net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11341__A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ net1321 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_10542_ net1 _06284_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13261_ net1320 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ team_03_WB.instance_to_wrap.wb.curr_state\[2\] team_03_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14149__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15000_ clknet_leaf_126_wb_clk_i net48 _01365_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12212_ net1596 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09766__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ net1351 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input68_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08650__A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12143_ net1655 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12074_ _06780_ net471 net445 net2019 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a22o_1
XANTENNA__11325__A0 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11025_ net656 _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11876__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09533__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15138__1519 vssd1 vssd1 vccd1 vccd1 _15138__1519/HI net1519 sky130_fd_sc_hd__conb_1
XFILLER_0_40_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08741__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__C net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12976_ net1431 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11235__B net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14715_ clknet_leaf_14_wb_clk_i _02479_ _01080_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11927_ _06625_ net2701 net374 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07432__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14646_ clknet_leaf_92_wb_clk_i _02410_ _01011_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\]
+ sky130_fd_sc_hd__dfstp_1
X_11858_ net272 net2668 net383 vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[28\] net309 net689 vssd1
+ vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11789_ net2670 _06469_ net332 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__mux2_1
X_14577_ clknet_leaf_93_wb_clk_i _02341_ _00942_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[931\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ net1273 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
XANTENNA__11800__A1 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ net1331 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09757__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XANTENNA__10906__A3 net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15129_ net1510 vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12108__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__A1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ net1121 _03888_ _03889_ _03891_ net1130 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__a311o_1
XFILLER_0_43_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06902_ net1014 net1012 net1015 vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07882_ net1103 team_03_WB.instance_to_wrap.core.register_file.registers_state\[47\]
+ net898 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__or3_1
XANTENNA__11129__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__A1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ team_03_WB.instance_to_wrap.WRITE_I vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09621_ net582 _05543_ _05544_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_91_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09552_ _05391_ _05395_ net563 vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08503_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08496__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09483_ _03641_ _04503_ net539 _05424_ _03639_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__o311a_1
XFILLER_0_52_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11860__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[826\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06954__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10984__B net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08365_ net1056 _04304_ _04305_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__or3_1
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout422_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__A0 _05881_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1164_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _03256_ _03257_ net806 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08296_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[24\]
+ net984 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07247_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07178_ net1106 _03117_ _03118_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10358__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09212__A2 _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08470__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout889_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11100__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07774__A2 net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1307 net1317 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout320 _05928_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_2
Xfanout1318 net1319 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_15_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1329 net1330 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__buf_4
XFILLER_0_10_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout331 _06811_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_6
XFILLER_0_22_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout353 net356 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12720__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 _06818_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_6
Xfanout375 net376 vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_8
XANTENNA__08184__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__buf_4
Xfanout397 net398 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_8
X_09819_ _02892_ net589 _04821_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12830_ net1414 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11055__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ net1355 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
X_14500_ clknet_leaf_19_wb_clk_i _02264_ _00865_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[854\]
+ sky130_fd_sc_hd__dfrtp_1
X_11712_ net2087 _06409_ net341 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
X_12692_ net1321 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10833__A2 _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12035__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14431_ clknet_leaf_114_wb_clk_i _02195_ _00796_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[785\]
+ sky130_fd_sc_hd__dfrtp_1
X_11643_ net1240 _06462_ net387 vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09987__A0 _05872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14362_ clknet_leaf_22_wb_clk_i _02126_ _00727_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _06447_ _06394_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08083__C net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
X_10525_ net1770 net1025 net1022 team_03_WB.instance_to_wrap.CPU_DAT_I\[14\] vssd1
+ vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ net1284 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
Xinput39 gpio_in[14] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14293_ clknet_leaf_90_wb_clk_i _02057_ _00658_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13244_ net1352 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
X_10456_ _06051_ _06052_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11546__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ net1416 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XANTENNA__11010__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] _06143_ vssd1 vssd1
+ vccd1 vccd1 _06215_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12126_ net1627 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14934__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08962__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _06623_ net2433 net363 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap318_A _05611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15113__1494 vssd1 vssd1 vccd1 vccd1 _15113__1494/HI net1494 sky130_fd_sc_hd__conb_1
XANTENNA__08714__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__A net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ net711 net701 net301 vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__or3b_1
XFILLER_0_75_1538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12959_ net1375 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13461__A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08573__S0 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14314__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10824__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__B1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14629_ clknet_leaf_124_wb_clk_i _02393_ _00994_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09978__A0 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08150_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\]
+ net949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\] net913
+ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10588__B2 _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07101_ net1140 _03042_ _03036_ net719 vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a211o_2
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07453__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08081_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[950\]
+ net892 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09386__A _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ net1183 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\]
+ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07205__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08402__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08983_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[10\] net995
+ net914 _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__o211a_1
XANTENNA__11855__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ net808 _03871_ _03872_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09053__S1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__C1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[443\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[315\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\]
+ net780 net1127 vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07064__S0 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07796_ _03733_ _03734_ net743 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _05371_ _05463_ _05468_ _05472_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_133_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout637_A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1379_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09466_ net550 _04417_ _05094_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08465__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08417_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\] net918
+ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09397_ _05170_ _05174_ _05338_ _05172_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[437\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[405\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[309\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[277\]
+ net959 net1067 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15137__1518 vssd1 vssd1 vccd1 vccd1 _15137__1518/HI net1518 sky130_fd_sc_hd__conb_1
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11240__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ net1213 _04220_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10310_ team_03_WB.instance_to_wrap.core.pc.current_pc\[29\] team_03_WB.instance_to_wrap.core.pc.current_pc\[28\]
+ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__A _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net506 net631 _06712_ net416 net2052 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a32o_1
XANTENNA__08619__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11528__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _06082_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07247__C net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1105 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06955__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1115 net1117 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__clkbuf_4
Xfanout1126 net1128 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_4
X_14980_ clknet_leaf_56_wb_clk_i _02732_ _01345_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dfrtp_1
Xfanout1137 team_03_WB.instance_to_wrap.core.ru.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net1137 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1148 net1150 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_4
Xfanout1159 net1160 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_4
XANTENNA__08157__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13931_ clknet_leaf_17_wb_clk_i _01695_ _00296_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07904__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14337__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ clknet_leaf_76_wb_clk_i _01626_ _00227_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[216\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12813_ net1318 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ clknet_leaf_1_wb_clk_i _01557_ _00158_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08555__S0 net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ net1351 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09614__A2_N _02803_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12675_ net1300 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14414_ clknet_leaf_68_wb_clk_i _02178_ _00779_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11626_ _06700_ net392 net355 net2644 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a22o_1
XANTENNA__11767__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ clknet_leaf_59_wb_clk_i _02109_ _00710_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09918__B _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08632__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ net656 _06667_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10508_ net2272 net1029 net1020 team_03_WB.instance_to_wrap.CPU_DAT_I\[31\] vssd1
+ vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a22o_1
Xhold609 team_03_WB.instance_to_wrap.core.register_file.registers_state\[258\] vssd1
+ vssd1 vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11488_ net1240 _06449_ net649 _06463_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__or4_4
X_14276_ clknet_leaf_12_wb_clk_i _02040_ _00641_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[630\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10990__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10439_ net284 _06137_ _06257_ net679 vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__o31ai_1
X_13227_ net1272 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10145__A _03109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13158_ net1423 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
XANTENNA__10742__A1 _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11675__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ net1134 net1137 team_03_WB.instance_to_wrap.core.ru.state\[5\] _06281_ net838
+ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__a221o_1
X_13089_ net1266 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08148__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11298__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08699__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09360__A1 _05278_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08163__A2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[654\] net760
+ net736 _03591_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07581_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[792\] net798
+ _02871_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11126__D net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09112__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09320_ _05259_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_111_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _05183_ _05187_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07674__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11470__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08202_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1011\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09182_ _03061_ _03062_ _03066_ _03104_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__and4b_1
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11758__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _03137_ _03170_ _04073_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nand4_4
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08064_ net1153 _04004_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__o21a_1
XANTENNA__11773__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07015_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\]
+ net876 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09179__B2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1127_A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__C1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08926__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09844__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__C1 _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07067__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11585__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13366__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ _04902_ _04907_ net869 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07917_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\] net782
+ _03858_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08897_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[236\] net935
+ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07848_ _03788_ _03789_ net609 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07779_ net807 _03719_ _03720_ net813 vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09103__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09518_ _05379_ _05382_ net563 vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10790_ _02829_ net688 _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07114__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11997__A0 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__C1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11333__B net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09449_ net547 net357 _05108_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o21ba_1
XANTENNA__07530__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ net1297 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11749__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15112__1493 vssd1 vssd1 vccd1 vccd1 _15112__1493/HI net1493 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _06468_ net2678 net401 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12391_ net1389 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08614__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11342_ net515 net635 _06723_ net408 net1843 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14130_ clknet_leaf_101_wb_clk_i _01894_ _00495_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07512__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10972__B2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11273_ net709 net298 net823 vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__and3_1
X_14061_ clknet_leaf_110_wb_clk_i _01825_ _00426_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13012_ net1322 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
X_10224_ _06012_ _06065_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
XANTENNA_input50_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11921__A0 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] net670 vssd1 vssd1 vccd1
+ vccd1 _05997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14963_ clknet_leaf_41_wb_clk_i _02715_ _01328_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__dfrtp_1
Xhold6 team_03_WB.instance_to_wrap.core.register_file.registers_state\[953\] vssd1
+ vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10086_ _05718_ _05730_ _05746_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10488__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ clknet_leaf_21_wb_clk_i _01678_ _00279_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14894_ clknet_leaf_44_wb_clk_i _02657_ _01259_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09893__A2 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ clknet_leaf_89_wb_clk_i _01609_ _00210_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11524__A _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13776_ clknet_leaf_83_wb_clk_i _01540_ _00141_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[130\]
+ sky130_fd_sc_hd__dfrtp_1
X_10988_ net2630 net427 _06565_ net506 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
XANTENNA__11988__A0 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11243__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12727_ net1415 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07656__A1 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08853__B1 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10660__A0 team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09929__A _03277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ net1403 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11609_ net649 net465 vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12589_ net1301 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08700__S0 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11755__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14328_ clknet_leaf_11_wb_clk_i _02092_ _00693_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold406 _02624_ vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold417 net198 vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\] vssd1
+ vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 net218 vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14259_ clknet_leaf_109_wb_clk_i _02023_ _00624_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08369__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09030__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout908 net909 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__clkbuf_4
Xfanout919 _04088_ vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08820_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\] net976
+ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__or2_1
XANTENNA__07041__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07592__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1106 team_03_WB.instance_to_wrap.core.register_file.registers_state\[783\] vssd1
+ vssd1 vccd1 vccd1 net2690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\] vssd1
+ vssd1 vccd1 vccd1 net2701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\] vssd1
+ vssd1 vccd1 vccd1 net2712 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _04687_ _04692_ net869 vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__mux2_1
XANTENNA__07615__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1139 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\] vssd1
+ vssd1 vccd1 vccd1 net2723 sky130_fd_sc_hd__dlygate4sd3_1
X_07702_ net1086 net891 team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\]
+ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__o21a_1
X_15136__1517 vssd1 vssd1 vccd1 vccd1 _15136__1517/HI net1517 sky130_fd_sc_hd__conb_1
X_08682_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[552\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__mux2_1
XANTENNA__07344__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07895__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\]
+ net788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\] net728
+ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11691__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07564_ _03504_ _03505_ net819 vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__o21a_1
XANTENNA__11979__A0 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09303_ _04591_ _05243_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__nor2_1
XANTENNA__07647__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07495_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[583\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\] net749
+ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout335_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1077_A _02788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09234_ _04235_ _05175_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ net577 _05106_ _05093_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09558__B _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout502_A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08116_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[858\]
+ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09096_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[877\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[845\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold940 team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\] vssd1
+ vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\] vssd1
+ vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[615\] vssd1
+ vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold973 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\] vssd1
+ vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold984 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[27\] vssd1 vssd1 vccd1
+ vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\] vssd1
+ vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11609__A net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _05883_ net2101 net288 vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08780__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ net869 _04889_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11960_ net621 _06737_ net461 net370 net2347 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a32o_1
XFILLER_0_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09875__A2 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ net313 net311 net321 _02780_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__a31o_1
XANTENNA__07886__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net634 _06700_ net472 net380 net2003 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13630_ net1400 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XANTENNA__09088__B1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10890__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _06442_ net2507 net521 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XANTENNA__08129__S net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09627__A2 _05568_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11063__B net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ net1426 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10773_ _02802_ _02807_ _02822_ _02827_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__or4_1
XFILLER_0_94_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10642__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ net1377 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XANTENNA_input98_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ net1334 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12443_ net1360 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07269__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15162_ net1543 vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_2
XANTENNA__08063__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ net1344 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08091__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ clknet_leaf_0_wb_clk_i _01877_ _00478_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07271__C1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ net265 net2842 net411 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__mux2_1
X_15093_ net1474 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
X_11256_ net501 net622 _06695_ net414 net2056 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a32o_1
X_14044_ clknet_leaf_128_wb_clk_i _01808_ _00409_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[398\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06901__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _06046_ _06048_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11187_ net508 net653 _06674_ net419 net1979 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11370__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10138_ _04119_ _02772_ net670 vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14946_ clknet_leaf_38_wb_clk_i _00008_ _01311_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10069_ _02825_ _05910_ _05911_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08523__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07877__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14877_ clknet_leaf_52_wb_clk_i _02640_ _01242_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13828_ clknet_leaf_12_wb_clk_i _01592_ _00193_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[182\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08266__C _04207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13759_ clknet_leaf_121_wb_clk_i _01523_ _00124_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11425__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10633__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07280_ _03218_ _03219_ net809 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11189__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08054__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 team_03_WB.instance_to_wrap.ADR_I\[23\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold214 _02591_ vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\] vssd1
+ vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 net221 vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 net230 vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold258 _02594_ vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _05435_ _05453_ _05500_ _05843_ _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__o2111ai_1
XANTENNA__07907__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__A _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold269 team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\] vssd1
+ vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09003__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout705 net708 vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__buf_4
Xfanout716 _06460_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
Xfanout727 net728 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
X_09852_ net579 _05683_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 net742 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__buf_4
XANTENNA__07565__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_4
X_08803_ net1046 team_03_WB.instance_to_wrap.core.register_file.registers_state\[65\]
+ net1000 team_03_WB.instance_to_wrap.core.register_file.registers_state\[97\] net939
+ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a221o_1
XANTENNA__11148__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__A3 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__C net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ _03459_ _04619_ _04816_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a21oi_1
X_06995_ _02925_ _02927_ _02932_ _02934_ _02926_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o2111a_4
XANTENNA_fanout285_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ net1214 _04672_ _04675_ net1073 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__o211a_1
X_15111__1492 vssd1 vssd1 vccd1 vccd1 _15111__1492/HI net1492 sky130_fd_sc_hd__conb_1
XFILLER_0_119_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10987__B net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07868__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _04601_ _04606_ net871 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout452_A _06801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11164__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07616_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\] net783
+ net749 _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a211o_1
XANTENNA__10872__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08596_ _02954_ _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07547_ _03460_ _03488_ net612 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux2_4
XANTENNA__08817__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1361_A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout717_A _02864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\] net762
+ net1037 vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11967__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09217_ _03567_ _03904_ _05155_ _02937_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_17_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11103__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07089__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08045__A1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ net439 net430 _04119_ net552 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__C1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ net858 _05017_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11110_ net830 net269 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__and2_2
XFILLER_0_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ _06789_ net481 net446 net2123 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold770 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\] vssd1
+ vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\] vssd1
+ vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net640 _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__nor2_1
XANTENNA__11339__A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[743\] vssd1
+ vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11352__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07556__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14800_ clknet_leaf_32_wb_clk_i _02564_ _01165_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07308__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ net1408 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10897__B _05821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07552__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ clknet_leaf_16_wb_clk_i _02495_ _01096_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11943_ net624 _06720_ net458 net369 net2799 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11074__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14662_ clknet_leaf_78_wb_clk_i _02426_ _01027_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11874_ net266 net2388 net383 vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13613_ net1281 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XANTENNA__08808__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[25\] net307 _06428_ net690
+ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__o211a_1
XFILLER_0_95_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14593_ clknet_leaf_1_wb_clk_i _02357_ _00958_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__D1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11958__A3 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ net1273 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
X_10756_ net2316 net532 net527 _06371_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12080__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11521__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13475_ net1399 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ _06314_ _06325_ net604 vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15214_ net910 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_1
X_12426_ net1256 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
XANTENNA__08036__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15135__1516 vssd1 vssd1 vccd1 vccd1 _15135__1516/HI net1516 sky130_fd_sc_hd__conb_1
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09784__A1 _03459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ net1526 vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
X_12357_ net1276 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09784__B2 _02945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11308_ _06618_ net2602 net412 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__mux2_1
X_15076_ net1457 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_121_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12288_ net1385 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
X_14027_ clknet_leaf_17_wb_clk_i _01791_ _00392_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A _03985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ net1242 net832 _06413_ net668 vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__and4_1
XANTENNA__07547__A0 _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08744__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14929_ clknet_leaf_125_wb_clk_i _02684_ _01294_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08450_ _04387_ _04388_ net855 vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07401_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[863\]
+ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08381_ net845 _04309_ _04322_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__o21a_4
XFILLER_0_4_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11134__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12808__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07332_ net1144 _03271_ _03272_ net1108 vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a31o_1
XANTENNA__11949__A3 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08275__A1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07263_ net723 _03188_ _03197_ _03204_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09002_ _04940_ _04943_ net1199 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11150__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ _03122_ _03135_ net720 vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_4
XFILLER_0_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11858__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09775__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07250__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09904_ _05844_ _05454_ _05429_ _05542_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__or4bb_2
XANTENNA__11159__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout502 net503 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
Xfanout524 _06395_ vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11334__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07538__B1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout535 net537 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout546 _03106_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__buf_2
X_09835_ _04566_ _04593_ net563 vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__o21a_1
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_2
XANTENNA__14220__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11593__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_A _06564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09571__B _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _05239_ _05271_ _05273_ net592 vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__a31o_1
X_06978_ net808 _02916_ _02918_ _02919_ net815 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__o311a_1
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08717_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[484\] net1073
+ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__a221o_1
XANTENNA__08189__S1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11637__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout834_A _06386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ _03866_ _05012_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09998__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10002__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08648_ _04582_ _04583_ _04589_ _04586_ net1061 net1077 vssd1 vssd1 vccd1 vccd1 _04590_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13938__CLK clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08579_ _04519_ _04520_ net1211 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10610_ net1621 team_03_WB.instance_to_wrap.CPU_DAT_O\[19\] net836 vssd1 vssd1 vccd1
+ vccd1 _02518_ sky130_fd_sc_hd__mux2_1
XANTENNA__09299__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08407__S net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _06477_ net2447 net452 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11341__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ net1684 net1030 net1021 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11270__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ net1299 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ team_03_WB.instance_to_wrap.wb.curr_state\[2\] team_03_WB.instance_to_wrap.wb.curr_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__nor2_2
XFILLER_0_106_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09215__B1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net1635 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13549__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ net1401 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11573__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12142_ net1623 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12073_ _05908_ _06394_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__nand2b_1
XANTENNA__08726__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ net1040 net834 net300 net669 vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14713__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07282__A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ net1388 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XANTENNA__11628__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14714_ clknet_leaf_118_wb_clk_i _02478_ _01079_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_11926_ _06624_ net2721 net374 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11235__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ clknet_leaf_72_wb_clk_i _02409_ _01010_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_129_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10847__S net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ _06681_ net466 net381 net2066 vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11532__A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[28\] net307 vssd1
+ vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__nand2_1
XANTENNA__08257__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14576_ clknet_leaf_80_wb_clk_i _02340_ _00941_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11788_ net2705 _06454_ net332 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
X_13527_ net1280 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XANTENNA__11251__B net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10739_ net2606 net531 net526 _06361_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09937__A _03563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ net1333 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
XANTENNA__07480__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15110__1491 vssd1 vssd1 vccd1 vccd1 _15110__1491/HI net1491 sky130_fd_sc_hd__conb_1
XANTENNA__09757__A1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ net1354 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
X_13389_ net1402 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_11_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11564__B2 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__07457__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15128_ net1509 vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
XFILLER_0_10_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
X_07950_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\]
+ net901 vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__or3_1
X_15059_ net1440 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XANTENNA__08717__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ net1016 net693 _02838_ _02841_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or4_4
X_07881_ _03821_ _03822_ net608 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_2
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11129__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _05549_ _05561_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2_2
X_06832_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] vssd1 vssd1 vccd1 vccd1
+ _02775_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14393__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07940__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _05392_ _05416_ net556 vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__mux2_1
XANTENNA__11619__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10827__A0 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08502_ _04430_ _04443_ net843 vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__mux2_4
XANTENNA__08496__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ _03641_ _04503_ net663 _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_A clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08433_ net1199 _04371_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or3_1
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08364_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\]
+ net960 net1067 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07315_ net1087 team_03_WB.instance_to_wrap.core.register_file.registers_state\[669\]
+ net727 _03245_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11252__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10055__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ net440 net429 _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout415_A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1157_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07246_ _03180_ _03187_ net1156 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__mux2_1
XANTENNA__07471__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11588__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\]
+ net756 net1116 vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1324_A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07759__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__A1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1308 net1309 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__buf_4
Xfanout310 _05846_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
Xfanout1319 net1335 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
Xfanout321 net322 vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
Xfanout332 net336 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_6
XFILLER_0_100_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout343 _06807_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__buf_8
Xfanout354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_8
Xfanout365 net366 vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08184__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout376 _06814_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_6
Xfanout387 net392 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_4
X_09818_ _02892_ net589 net665 _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__a22o_1
Xfanout398 _06757_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_55_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10530__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _04775_ _05570_ net359 vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__o21bai_1
X_15134__1515 vssd1 vssd1 vccd1 vccd1 _15134__1515/HI net1515 sky130_fd_sc_hd__conb_1
XFILLER_0_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12760_ net1369 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XANTENNA__11055__C net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__B1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__S _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11711_ net1943 net281 net342 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ net1265 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14430_ clknet_leaf_57_wb_clk_i _02194_ _00795_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\]
+ sky130_fd_sc_hd__dfrtp_1
X_11642_ _06716_ net390 net355 net2455 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ clknet_leaf_103_wb_clk_i _02125_ _00726_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11573_ net2230 net489 _06799_ net516 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07998__B1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_1
XANTENNA__11794__A1 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input80_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ net1288 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
X_10524_ net2290 net1030 net1021 net1974 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14292_ clknet_leaf_92_wb_clk_i _02056_ _00657_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09739__A1 _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ net1360 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
XANTENNA__09739__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ net2874 _06270_ net679 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08411__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ net1338 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10386_ net2009 _06214_ net677 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07845__S0 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ net1631 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06973__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1443 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12056_ _06622_ net2736 net364 vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__mux2_1
XANTENNA__08600__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__C net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08175__B1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ net2628 net427 _06576_ net499 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XANTENNA__07216__S net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10809__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08478__A1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ net1386 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XANTENNA__08836__A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__B1 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08573__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11909_ _06609_ net2634 net376 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__mux2_1
XANTENNA__07150__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__A3 net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ net1355 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_14628_ clknet_leaf_16_wb_clk_i _02392_ _00993_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12026__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14609__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07438__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ clknet_leaf_114_wb_clk_i _02323_ _00924_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07100_ _03039_ _03040_ _03041_ net1110 vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08080_ _04019_ _04021_ net1153 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07031_ net1140 _02961_ _02972_ net718 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__a211oi_2
XANTENNA__13189__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11201__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08938__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14759__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08402__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07610__C1 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\] net954
+ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09606__S net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07933_ net743 _03873_ _03874_ net805 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08166__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ net814 _03804_ _03805_ _03797_ _03800_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a32o_1
XANTENNA__07064__S1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ _04828_ _05460_ net575 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__mux2_2
X_07795_ _03735_ _03736_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout365_A net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09115__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14139__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _04536_ _04777_ _05475_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09465_ _05405_ _05406_ net555 vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__A1 net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1274_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ net933 _04356_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__o21a_1
XANTENNA__12017__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _05331_ _05335_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07692__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14289__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08347_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\]
+ net959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\] net1202
+ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10579__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07796__S net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08278_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[407\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[311\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\]
+ net970 net1070 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout999_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07229_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__or3_1
XFILLER_0_127_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11528__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11111__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _03944_ _05998_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10171_ _06010_ _06011_ _03758_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06955__A1 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1105 _02787_ vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__clkbuf_4
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
XANTENNA__07825__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1127 net1128 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1138 net1141 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_6
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
XANTENNA__08157__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ clknet_leaf_9_wb_clk_i _01694_ _00295_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11347__A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13861_ clknet_leaf_106_wb_clk_i _01625_ _00226_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11066__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11781__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12812_ net1305 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ clknet_leaf_132_wb_clk_i _01556_ _00157_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12743_ net1398 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XANTENNA__08555__S1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__C1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07132__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11082__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12008__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ net1348 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11216__A0 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14413_ clknet_leaf_104_wb_clk_i _02177_ _00778_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[767\]
+ sky130_fd_sc_hd__dfrtp_1
X_11625_ _06699_ net388 net355 net2440 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13656__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ clknet_leaf_27_wb_clk_i _02108_ _00709_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07435__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ net497 net620 _06666_ net486 net1947 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__a32o_1
XANTENNA__08632__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08391__A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10507_ team_03_WB.instance_to_wrap.wb.curr_state\[1\] _02797_ team_03_WB.instance_to_wrap.wb.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3b_1
X_14275_ clknet_leaf_25_wb_clk_i _02039_ _00640_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[629\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11487_ net2624 net400 _06777_ net519 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
Xmax_cap318 _05611_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10990__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13226_ net1250 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
X_10438_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] _06136_ vssd1 vssd1 vccd1
+ vccd1 _06257_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ net1272 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
X_10369_ net286 _06146_ _06197_ net677 vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__o31a_1
XANTENNA__06946__B2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ net1137 net604 _06300_ net1687 net1134 vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a32o_1
XANTENNA__08330__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13088_ net1409 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11257__A _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _06777_ net483 net368 net2794 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08699__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09360__A2 _05281_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07371__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[28\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07580_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[824\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07470__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11455__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07123__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15205__1575 vssd1 vssd1 vccd1 vccd1 _15205__1575/HI net1575 sky130_fd_sc_hd__conb_1
XFILLER_0_34_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07123__B2 net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09250_ _05190_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11207__A0 _06438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08201_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[947\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\]
+ net948 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ net554 _04807_ _05121_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12816__A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14581__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08132_ _03208_ _03243_ _03759_ _03790_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__and4b_2
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08623__A1 net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08063_ net1118 _04000_ _04001_ _04003_ net1108 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15133__1514 vssd1 vssd1 vccd1 vccd1 _15133__1514/HI net1514 sky130_fd_sc_hd__conb_1
XFILLER_0_101_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09179__A2 _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07014_ net1182 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\]
+ net876 _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__A2 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ net1215 _04905_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout482_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11167__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07916_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[943\]
+ net881 _02870_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08896_ _04836_ _04837_ net857 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09860__A _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] net821 vssd1 vssd1 vccd1
+ vccd1 _03789_ sky130_fd_sc_hd__nand2_1
XANTENNA__11694__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1391_A net1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout747_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07778_ net726 _03708_ _03709_ _03707_ net802 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a311o_1
XANTENNA__07380__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ net563 _05380_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11106__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10010__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09448_ net591 _05340_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11333__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14924__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07665__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ _05315_ _05320_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11749__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ _06453_ net2585 net401 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ net1411 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08614__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ net303 net713 net699 vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ clknet_leaf_8_wb_clk_i _01824_ _00425_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\]
+ sky130_fd_sc_hd__dfrtp_1
X_11272_ net502 net621 _06703_ net414 net2149 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ net1259 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
X_10223_ _06017_ _06021_ _06062_ _06016_ _06013_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a311o_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_70_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_input43_A gpio_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14962_ clknet_leaf_31_wb_clk_i _02714_ _01327_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold7 team_03_WB.instance_to_wrap.core.register_file.registers_state\[936\] vssd1
+ vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
X_10085_ _05757_ _05926_ net321 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07889__C1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11685__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13913_ clknet_leaf_111_wb_clk_i _01677_ _00278_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14454__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14893_ clknet_leaf_43_wb_clk_i _02656_ _01258_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13844_ clknet_leaf_90_wb_clk_i _01608_ _00209_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[198\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07290__A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13775_ clknet_leaf_100_wb_clk_i _01539_ _00140_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10987_ net281 net653 net705 net826 vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ net1346 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XANTENNA__11243__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08853__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12657_ net1315 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11608_ net656 net472 vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12588_ net1298 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09010__A net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10412__A1 _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14327_ clknet_leaf_86_wb_clk_i _02091_ _00692_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08700__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ net2315 net487 _06787_ net505 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold407 net236 vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold418 team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\] vssd1
+ vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09945__A _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14258_ clknet_leaf_105_wb_clk_i _02022_ _00623_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold429 team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\] vssd1
+ vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08369__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13209_ net1357 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ clknet_leaf_106_wb_clk_i _01953_ _00554_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[543\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout909 _05906_ vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07041__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1107 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\] vssd1
+ vssd1 vccd1 vccd1 net2691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08750_ net1060 _04690_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1118 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\] vssd1
+ vssd1 vccd1 vccd1 net2702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\] vssd1
+ vssd1 vccd1 vccd1 net2713 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10479__B2 team_03_WB.instance_to_wrap.ADR_I\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08681_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\]
+ net978 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07632_ net1168 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\]
+ net873 _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__a31o_1
XANTENNA__13821__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11428__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ net1126 _03501_ _03502_ net1112 vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_113_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _04591_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07494_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[647\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ _03904_ _05156_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10651__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11450__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ net565 _05105_ _05100_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08115_ _04050_ _04051_ _04056_ net1154 vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o22a_1
XANTENNA__11600__A0 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09095_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1005\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[973\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__mux2_1
XANTENNA__10066__A team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1237_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07280__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08046_ _03986_ _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nor2_1
Xhold930 team_03_WB.instance_to_wrap.core.register_file.registers_state\[794\] vssd1
+ vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\] vssd1
+ vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11596__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\] vssd1
+ vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold963 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1 net2547
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09021__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1404_A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\] vssd1
+ vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11903__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\] vssd1
+ vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap693 _02834_ vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_1
Xhold996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\] vssd1
+ vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14477__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11609__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _05882_ net1966 net290 vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__mux2_1
XANTENNA__07583__A1 net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08780__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10005__S net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net921 _04887_ _04888_ net859 vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10910_ net691 _05676_ net586 vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__o21ai_1
X_11890_ net628 _06699_ net466 net378 net2022 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11419__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10890__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ _06439_ _06440_ _06441_ net586 vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__o211a_2
XFILLER_0_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ net1313 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XANTENNA__12092__B1 net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] net1240 vssd1 vssd1 vccd1
+ vccd1 _06382_ sky130_fd_sc_hd__nand2_1
XANTENNA__08934__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ net1374 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13491_ net1334 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08653__B net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ net1371 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ net1542 vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_2
XFILLER_0_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ net1262 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14112_ clknet_leaf_134_wb_clk_i _01876_ _00477_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11324_ _06629_ net2504 net411 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15092_ net1473 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14043_ clknet_leaf_34_wb_clk_i _01807_ _00408_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\]
+ sky130_fd_sc_hd__dfrtp_1
X_11255_ net274 net709 net822 vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ _04739_ net672 _06044_ _02994_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__o211ai_1
XANTENNA__07285__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ net705 _06532_ net699 vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _03528_ _05978_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14945_ clknet_leaf_38_wb_clk_i _00007_ _01310_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10068_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] team_03_WB.instance_to_wrap.core.decoder.inst\[13\]
+ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] team_03_WB.instance_to_wrap.core.decoder.inst\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08523__B1 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09866__A3 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14876_ clknet_leaf_50_wb_clk_i _02639_ _01241_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15132__1513 vssd1 vssd1 vccd1 vccd1 _15132__1513/HI net1513 sky130_fd_sc_hd__conb_1
XANTENNA__09079__A1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07451__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ clknet_leaf_19_wb_clk_i _01591_ _00192_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13758_ clknet_leaf_48_wb_clk_i _01522_ _00123_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08826__A1 net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08844__A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10633__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12709_ net1276 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11830__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13689_ clknet_leaf_83_wb_clk_i _01453_ _00054_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11189__A2 net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold204 _02626_ vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold215 team_03_WB.instance_to_wrap.core.register_file.registers_state\[52\] vssd1
+ vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07262__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 net214 vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\] vssd1
+ vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold248 net212 vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ _05847_ _05596_ _05583_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__nor3b_1
Xhold259 team_03_WB.instance_to_wrap.core.register_file.registers_state\[699\] vssd1
+ vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09003__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_4
X_09851_ net564 _05136_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__nor2_1
XANTENNA__08211__C1 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout717 _02864_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__clkbuf_8
Xfanout728 net736 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
XANTENNA__11897__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07626__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout739 net741 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
X_08802_ _04742_ _04743_ net852 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__o21a_1
X_09782_ net580 _05638_ _05723_ net360 vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__o211a_1
XANTENNA__11148__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06994_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] _02832_ _02925_ _02927_
+ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__nor4_1
XANTENNA__07923__A _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[868\] net1061
+ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__C net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08664_ net1062 _04604_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07615_ net1195 team_03_WB.instance_to_wrap.core.register_file.registers_state\[569\]
+ net881 vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and3_1
XANTENNA__11164__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10872__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08595_ _04327_ _04536_ net581 vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1187_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12074__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07546_ net718 _03471_ _03480_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o22a_4
XFILLER_0_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08817__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07477_ _03417_ _03418_ net1154 vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07096__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1092 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1354_A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ net605 _03529_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ _05087_ _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__S0 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__A2 _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07253__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ net851 _05018_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08029_ net742 _03969_ _03970_ _02849_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a31o_1
Xhold760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\] vssd1
+ vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\] vssd1
+ vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold782 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\] vssd1
+ vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11040_ net702 net713 net297 vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__or3b_1
Xhold793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\] vssd1
+ vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__B net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07556__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11352__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10560__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12991_ net1377 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XANTENNA__07308__A1 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__A _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14730_ clknet_leaf_42_wb_clk_i _02494_ _01095_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ net631 _06719_ net471 net372 net2403 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11074__B net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14661_ clknet_leaf_124_wb_clk_i _02425_ _01026_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\]
+ sky130_fd_sc_hd__dfstp_1
X_11873_ net267 net2232 net382 vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ net1273 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10824_ net313 net311 net322 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a31o_1
X_14592_ clknet_leaf_133_wb_clk_i _02356_ _00957_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08808__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10076__C1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13543_ net1327 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] _05757_ net603 vssd1
+ vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__mux2_1
XANTENNA__11812__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13474_ net1399 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10686_ _06319_ _06326_ net600 vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__a21o_1
X_15213_ net1578 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12425_ net1252 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ net1525 vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
XFILLER_0_50_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07244__B1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ net1306 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09784__A2 _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06912__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08603__S net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11307_ _06617_ net2683 net412 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15075_ net1456 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
X_12287_ net1374 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XANTENNA__14792__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14026_ clknet_leaf_4_wb_clk_i _01790_ _00391_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ net496 net617 _06686_ net413 net2402 vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a32o_1
XANTENNA__11879__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A1 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08744__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11169_ net2576 net418 _06663_ net501 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
XANTENNA__11894__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14928_ clknet_leaf_39_wb_clk_i _02683_ _01293_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14859_ clknet_leaf_54_wb_clk_i net1732 _01224_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13480__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__A0 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[895\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08380_ net863 _04321_ _04316_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08574__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07331_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\]
+ net767 net1120 vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07262_ net814 _03203_ net719 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ net1208 _04941_ _04942_ net1066 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07193_ net1138 _03129_ _03134_ net812 vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09775__A2 _05485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__B2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08432__C1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08983__B1 net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07786__B2 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10790__B1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ _05844_ _05455_ _05429_ _05542_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11159__B net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout514 _06448_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
Xfanout525 net528 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11874__S net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08735__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11334__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 net549 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
X_09834_ net327 _05436_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_127_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout558 net560 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06968__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08749__A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout569 _03025_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
X_09765_ _05239_ _05271_ _05273_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__a21oi_1
X_06977_ _02914_ _02915_ net805 vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11175__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08716_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\] net1204
+ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a221o_1
X_09696_ _04150_ _04326_ _05014_ _04210_ net561 net574 vssd1 vssd1 vccd1 vccd1 _05638_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08647_ _04587_ _04588_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__A1 net1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07171__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08578_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\]
+ net965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\] net933
+ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14665__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07529_ _03463_ _03464_ _03469_ _03470_ net1110 net1131 vssd1 vssd1 vccd1 vccd1 _03471_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11114__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ net171 net1024 net905 net1585 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
XANTENNA__07474__B1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11270__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08671__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10471_ net1135 net2104 _06282_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__o21a_1
XANTENNA__12734__A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ net1594 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ net1423 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XANTENNA__07777__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11573__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net1674 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__clkbuf_1
X_15131__1512 vssd1 vssd1 vccd1 vccd1 _15131__1512/HI net1512 sky130_fd_sc_hd__conb_1
XFILLER_0_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14045__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ _06633_ net2537 net363 vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold590 team_03_WB.instance_to_wrap.core.register_file.registers_state\[283\] vssd1
+ vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11784__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ net515 net658 _06585_ net427 net1937 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10533__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11876__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14195__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ net1337 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1290 team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] vssd1 vssd1 vccd1 vccd1
+ net2874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713_ clknet_leaf_11_wb_clk_i _02477_ _01078_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_11925_ _06623_ net2747 net375 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07162__C1 _02843_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12909__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11856_ net273 net2217 net381 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__mux2_1
X_14644_ clknet_leaf_91_wb_clk_i _02408_ _01009_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[998\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06907__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10807_ _06413_ net2765 net521 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__mux2_1
X_14575_ clknet_leaf_98_wb_clk_i _02339_ _00940_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[929\]
+ sky130_fd_sc_hd__dfrtp_1
X_11787_ net2502 _06620_ net332 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10738_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] _05697_ net603 vssd1
+ vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07465__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13526_ net1281 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XANTENNA__11251__C net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13457_ net1331 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09206__A1 _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09937__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ _05455_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12408_ net1362 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XANTENNA__09757__A2 _04922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07738__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ net1400 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XANTENNA__08333__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XANTENNA__11564__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
X_15127_ net1508 vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_2
XFILLER_0_2_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12339_ net1261 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XANTENNA__10164__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09953__A _03984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15058_ net1439 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__08717__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14009_ clknet_leaf_103_wb_clk_i _01773_ _00374_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\]
+ sky130_fd_sc_hd__dfrtp_1
X_06900_ net1016 net693 _02838_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nor4_2
XFILLER_0_120_1450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07880_ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] net1017 net682 vssd1
+ vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10524__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14538__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__A net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08193__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06831_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] vssd1 vssd1 vccd1 vccd1
+ _02774_ sky130_fd_sc_hd__inv_2
X_09550_ _03529_ _04267_ net539 _05491_ _03527_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__o311a_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09142__A0 _04149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08501_ _04437_ _04442_ net869 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09481_ _03641_ _04503_ net541 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07153__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08432_ net933 _04373_ _04372_ net1056 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12029__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\] net1202
+ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__o221a_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07314_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\] net767
+ net740 _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__a211o_1
XANTENNA__11252__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08294_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11869__S net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ net1131 _03181_ _03182_ _03185_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout310_A _05846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12554__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11004__B2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07176_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\]
+ net754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o221a_1
XANTENNA__14068__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07759__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11555__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1317_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout300 _06487_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
Xfanout311 net312 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_4
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout777_A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout322 net323 vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout333 net335 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_6
XANTENNA__10515__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08184__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 net356 vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_6
XFILLER_0_103_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout366 _06817_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_4
Xfanout377 net378 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_8
X_09817_ net584 net589 net543 vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13905__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout388 net392 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_4
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__S net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ net585 _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ _05568_ _05514_ _05355_ _05565_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11055__D net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11710_ _06459_ _06803_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__or2_4
XFILLER_0_96_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ net1398 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07695__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07790__S0 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ _06715_ net389 net354 net2409 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12035__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ clknet_leaf_8_wb_clk_i _02124_ _00725_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\]
+ sky130_fd_sc_hd__dfrtp_1
X_11572_ net642 net708 net266 net698 vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11779__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__S0 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ net1293 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
X_10523_ net143 net1030 net1021 net1780 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
X_14291_ clknet_leaf_109_wb_clk_i _02055_ _00656_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13242_ net1365 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XANTENNA_input73_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ net284 _06054_ _06269_ _06268_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a31o_1
XANTENNA__09739__A2 _04953_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__B1 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13173_ net1269 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
X_10385_ _06211_ _06213_ net283 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07845__S1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12124_ net1698 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09773__A net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12055_ _06479_ net2525 net362 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09923__D _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net653 _06575_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__and2_1
XANTENNA__07293__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07922__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[28\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09675__A1 _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ net1382 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__B2 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11908_ net1040 net653 _06463_ net468 vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__or4b_4
XANTENNA__07686__B1 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__B _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08328__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12888_ net1369 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14627_ clknet_leaf_25_wb_clk_i _02391_ _00992_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10159__A _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ net655 _06677_ net469 net329 net1880 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a32o_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10037__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07438__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ clknet_leaf_57_wb_clk_i _02322_ _00923_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13509_ net1325 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14489_ clknet_leaf_111_wb_clk_i _02253_ _00854_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07030_ _02963_ _02966_ _02971_ net1110 net1131 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__o221a_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11537__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09060__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ net443 net435 _04922_ net554 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__o31a_1
X_07932_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\]
+ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08166__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ net804 _03793_ _03794_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__or3_1
XFILLER_0_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09602_ _05171_ _05172_ _05174_ _05338_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o211ai_2
X_07794_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\] net730
+ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__a221o_1
XANTENNA__09115__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ _03566_ _04354_ net539 _05474_ _03564_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__o311a_1
XANTENNA__07931__A net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09666__B2 net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout358_A _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ net550 _04384_ _05096_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__a21oi_1
X_15130__1511 vssd1 vssd1 vccd1 vccd1 _15130__1511/HI net1511 sky130_fd_sc_hd__conb_1
XANTENNA__07141__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[186\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[154\] net961 net919
+ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09395_ _05174_ _05336_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout525_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08346_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\]
+ net959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[373\] net1067
+ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__o221a_1
XANTENNA__07429__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11225__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11599__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[471\]
+ net969 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14703__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07228_ _03139_ _03169_ net610 vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__mux2_2
XFILLER_0_105_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout894_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08929__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11528__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10008__S net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ net819 _03096_ _03098_ _03100_ net722 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__a41o_1
XFILLER_0_28_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09051__C1 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10170_ _03758_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1117 _02785_ vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
XANTENNA__08157__A1 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__clkbuf_4
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_4
XANTENNA__11347__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__A _03943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A2 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ clknet_leaf_8_wb_clk_i _01624_ _00225_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[214\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09106__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12811_ net1271 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ clknet_leaf_121_wb_clk_i _01555_ _00156_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12110__C1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07668__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12742_ net1419 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11082__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12673_ net1288 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08880__A2 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ _06698_ net385 net353 net2326 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
X_14412_ clknet_leaf_7_wb_clk_i _02176_ _00777_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08617__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11767__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14343_ clknet_leaf_68_wb_clk_i _02107_ _00708_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\]
+ sky130_fd_sc_hd__dfrtp_1
X_11555_ net2233 net488 _06792_ net508 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11302__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__B net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ net1965 net1027 net903 net1896 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_745 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14274_ clknet_leaf_131_wb_clk_i _02038_ _00639_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\]
+ sky130_fd_sc_hd__dfrtp_1
X_11486_ net642 net707 net266 net826 vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ net1247 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
X_10437_ _06057_ _06059_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10727__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12922__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13156_ net1307 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
X_10368_ net305 net304 _06198_ _06199_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ _02765_ net1739 _06820_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11538__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13087_ net1378 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
X_10299_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] _06140_ vssd1 vssd1
+ vccd1 vccd1 _06141_ sky130_fd_sc_hd__and2_1
XANTENNA__08148__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__B2 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ _06776_ net478 net367 net2399 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__a22o_1
XANTENNA__11257__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07356__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07751__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07108__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13989_ clknet_leaf_108_wb_clk_i _01753_ _00354_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11273__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08200_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09180_ net553 _04807_ net540 net665 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o31ai_1
XANTENNA__14726__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__A2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _03604_ _03728_ _03866_ _03990_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__and4b_1
XANTENNA__08084__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11212__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08062_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[406\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[278\]
+ net766 net1119 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14876__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07013_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\]
+ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09033__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08387__A1 net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__B2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A1 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11448__A _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12043__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ net1063 _04903_ _04904_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07915_ _03854_ _03856_ net1112 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__a21o_1
XANTENNA__11167__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[172\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\] net958 net917
+ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a221o_1
XANTENNA__10071__B _05914_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout475_A net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10497__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07846_ net717 _03787_ _03776_ _03768_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_58_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07661__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ net739 _03716_ _03717_ _03718_ _03702_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout642_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1384_A net1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ net558 _05375_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08847__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08311__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _05167_ _05339_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout907_A _05907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09378_ _05318_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[757\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[725\]
+ net962 vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10957__B1 net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ net497 net618 _06722_ net405 net2318 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a32o_1
XANTENNA__07822__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09024__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ net709 net299 net822 vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13010_ net1420 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10222_ _06016_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08431__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _03985_ _05993_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14961_ clknet_leaf_31_wb_clk_i _02713_ _01326_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__dfrtp_1
XANTENNA_input36_A gpio_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _05082_ _05142_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09878__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__S net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_03_WB.instance_to_wrap.core.register_file.registers_state\[982\] vssd1
+ vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13912_ clknet_leaf_118_wb_clk_i _01676_ _00277_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07889__B1 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ clknet_leaf_43_wb_clk_i _02655_ _01257_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13843_ clknet_leaf_112_wb_clk_i _01607_ _00208_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11093__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__B2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14749__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10986_ _06463_ net694 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__nand2_2
XANTENNA__11524__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13774_ clknet_leaf_71_wb_clk_i _01538_ _00139_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[128\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12725_ net1260 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12656_ net1427 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XANTENNA__08606__S net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14899__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13773__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ _06557_ net2643 net455 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12587_ net1257 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09802__A1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10412__A2 _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07813__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14326_ clknet_leaf_84_wb_clk_i _02090_ _00691_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11538_ net652 _06648_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold408 team_03_WB.instance_to_wrap.core.register_file.registers_state\[438\] vssd1
+ vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold419 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\] vssd1
+ vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ clknet_leaf_96_wb_clk_i _02021_ _00622_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[611\]
+ sky130_fd_sc_hd__dfrtp_1
X_11469_ net2663 net399 _06770_ net510 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08369__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13208_ net1368 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ clknet_leaf_8_wb_clk_i _01952_ _00553_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07041__A1 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13139_ net1264 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
Xhold1108 team_03_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1 net2692
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09869__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1119 team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\] vssd1
+ vssd1 vccd1 vccd1 net2703 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ net1086 net891 team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08680_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[680\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\]
+ net977 vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11046__C_N net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08541__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\]
+ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07895__A3 net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11207__S net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ net1158 _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09301_ _03489_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07493_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[551\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _04415_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08516__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09201__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09163_ _05102_ _05104_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08057__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ net740 _04052_ _04053_ _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[941\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XANTENNA__07804__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10066__B team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08045_ net717 _03962_ _03983_ net610 vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__o211a_1
XANTENNA__09006__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__A net1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold920 team_03_WB.instance_to_wrap.core.register_file.registers_state\[711\] vssd1
+ vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1132_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 team_03_WB.instance_to_wrap.core.register_file.registers_state\[809\] vssd1
+ vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold942 team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\] vssd1
+ vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold953 team_03_WB.instance_to_wrap.core.register_file.registers_state\[64\] vssd1
+ vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08251__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold964 team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\] vssd1
+ vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11364__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\] vssd1
+ vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold986 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\] vssd1
+ vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11178__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[397\] vssd1
+ vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10082__A _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _05881_ net2023 net288 vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__mux2_1
XANTENNA__08780__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08947_ _04885_ _04886_ net852 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11667__A1 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08878_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__and2b_4
XFILLER_0_135_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07829_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[458\]
+ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11117__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ net686 _05842_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10890__A2 _05646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__D_N _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10771_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] net1015 vssd1 vssd1 vccd1
+ vccd1 _06381_ sky130_fd_sc_hd__nand2_1
X_12510_ net1385 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
X_13490_ net1334 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08426__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09111__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12441_ net1356 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15160_ net1541 vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_2
X_12372_ net1322 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08950__A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11787__S net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14111_ clknet_leaf_115_wb_clk_i _01875_ _00476_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[465\]
+ sky130_fd_sc_hd__dfrtp_1
X_11323_ _06519_ net2390 net411 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__mux2_1
XANTENNA__07271__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15091_ net1472 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09548__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14042_ clknet_leaf_19_wb_clk_i _01806_ _00407_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ net504 net624 _06694_ net413 net2271 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a32o_1
XANTENNA__08161__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14421__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _05953_ _05956_ _05952_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11088__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11185_ net2183 net419 _06673_ net512 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10136_ _04267_ _02771_ net671 vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__A _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10067_ net1200 net1203 net1212 net1043 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__or4_1
X_14944_ clknet_leaf_124_wb_clk_i _02699_ _01309_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11658__A1 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14571__CLK clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08523__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14875_ clknet_leaf_52_wb_clk_i _02638_ _01240_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ clknet_leaf_131_wb_clk_i _01590_ _00191_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[180\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ clknet_leaf_68_wb_clk_i _01521_ _00122_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10969_ net690 _05082_ _06399_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ net1306 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XANTENNA__08336__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13688_ clknet_leaf_11_wb_clk_i _01452_ _00053_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08563__C _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ net1375 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11189__A3 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11594__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold205 team_03_WB.instance_to_wrap.ADR_I\[13\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13478__A net1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14309_ clknet_leaf_107_wb_clk_i _02073_ _00674_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[663\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07262__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold216 net197 vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 net185 vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold238 net205 vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 team_03_WB.instance_to_wrap.core.register_file.registers_state\[424\] vssd1
+ vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11346__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07907__C net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07014__A1 net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ net557 _05133_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nor2_1
XANTENNA__13669__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11897__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout729 net735 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[129\]
+ net975 team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\] net939
+ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__o221a_1
X_09781_ _02992_ _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or2_1
X_06993_ _02792_ _02927_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08732_ net1214 _04671_ _04673_ net1204 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__o211a_1
XANTENNA__09711__B1 _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10987__D net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ net1215 _04602_ _04603_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07614_ net1149 _03554_ _03555_ net819 vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__o31a_1
X_08594_ _04386_ _04448_ _04534_ _04478_ net564 net568 vssd1 vssd1 vccd1 vccd1 _04536_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10872__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ net818 _03486_ net723 vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1082_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_A _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07476_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[981\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1013\] net1143
+ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o221a_1
XFILLER_0_14_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11821__A1 net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ _03904_ _05155_ _02937_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__o21a_1
XFILLER_0_63_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1347_A net1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ net438 net430 _04236_ net544 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__o31a_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11585__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14444__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08676__S1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07253__A1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[205\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\] net933
+ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08450__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11400__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\]
+ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__or2_1
Xhold750 team_03_WB.instance_to_wrap.core.register_file.registers_state\[365\] vssd1
+ vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout974_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 team_03_WB.instance_to_wrap.ADR_I\[25\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\] vssd1
+ vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\] vssd1
+ vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\] vssd1
+ vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14594__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__C net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09979_ _03059_ net2138 net293 vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12990_ net1386 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
XANTENNA__11355__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11941_ _02793_ net658 _06562_ net472 vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or4b_4
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14660_ clknet_leaf_17_wb_clk_i _02424_ _01025_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1014\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ _06545_ net2193 net382 vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__mux2_1
XANTENNA__09540__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13611_ net1331 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10823_ net692 _05479_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ clknet_leaf_114_wb_clk_i _02355_ _00956_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[945\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_3_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11371__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08364__S0 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ net1273 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10754_ net527 _06369_ _06370_ net532 net1920 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09481__A2 _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10685_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] _06318_ vssd1 vssd1
+ vccd1 vccd1 _06326_ sky130_fd_sc_hd__or2_1
X_13473_ net1324 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15212_ net911 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07995__S net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12424_ net1285 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11576__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__A3 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15143_ net1524 vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
XFILLER_0_45_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07244__A1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12355_ net1296 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11310__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13811__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _06616_ net2625 net411 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__mux2_1
XANTENNA__11328__A0 _06631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15074_ net1455 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
X_12286_ net1384 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14025_ clknet_leaf_59_wb_clk_i _01789_ _00390_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[379\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237_ net280 net710 net822 vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11879__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__A0 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08744__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ net622 _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07952__C1 net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ _04504_ team_03_WB.instance_to_wrap.core.pc.current_pc\[30\] net671 vssd1
+ vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ net828 net298 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11265__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14927_ clknet_leaf_126_wb_clk_i _02682_ _01292_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11500__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11980__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14317__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14858_ clknet_leaf_41_wb_clk_i _02622_ _01223_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13809_ clknet_leaf_95_wb_clk_i _01573_ _00174_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14789_ clknet_leaf_41_wb_clk_i _02553_ _01154_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07330_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\]
+ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__or2_1
XANTENNA__11281__A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__A1 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07261_ net1156 _03201_ _03202_ _03200_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09000_ net1041 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\]
+ net994 team_03_WB.instance_to_wrap.core.register_file.registers_state\[874\] net1057
+ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07192_ _03130_ _03131_ _03132_ _03133_ net806 net724 vssd1 vssd1 vccd1 vccd1 _03134_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11031__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13001__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07786__A2 _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10790__A1 _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _05563_ _05824_ _05843_ _05583_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11159__C net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 net520 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_4
Xfanout526 net528 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
X_09833_ net592 _05771_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__o21ai_1
Xfanout548 net549 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout290_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 net560 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07943__C1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net592 _05698_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__o21a_2
X_06976_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\] net771
+ net729 _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08715_ net860 _04655_ _04656_ _04654_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__a31o_1
XANTENNA__11175__B net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09695_ _05196_ _05635_ _05203_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1297_A net1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__S0 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\] net922
+ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08577_ net1227 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\]
+ net966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[637\] net919
+ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _03465_ _03466_ net750 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ net806 _03396_ _03397_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11270__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ net1134 team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _06282_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08704__S _04097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07226__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09129_ _05042_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12140_ net1683 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12071_ _06632_ net2616 net363 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\] vssd1
+ vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 team_03_WB.instance_to_wrap.core.register_file.registers_state\[549\] vssd1
+ vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ net708 net272 net826 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__and3_1
XANTENNA__08726__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12973_ net1301 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1280 team_03_WB.instance_to_wrap.core.register_file.registers_state\[648\] vssd1
+ vssd1 vccd1 vccd1 net2864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1291 team_03_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1 net2875
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14712_ clknet_leaf_120_wb_clk_i _02476_ _01077_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ _06622_ net2413 net376 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14643_ clknet_leaf_115_wb_clk_i _02407_ _01008_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\]
+ sky130_fd_sc_hd__dfstp_1
X_11855_ _06468_ net2320 net381 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11305__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06907__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__S0 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10806_ _06410_ _06411_ _06412_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__a21o_1
XANTENNA__11532__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14574_ clknet_leaf_70_wb_clk_i _02338_ _00939_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\]
+ sky130_fd_sc_hd__dfrtp_1
X_11786_ net2458 _06619_ net332 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13525_ net1273 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10737_ net1789 net531 net525 _06360_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11251__D net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ net1332 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10668_ _05541_ _05932_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__nor2_1
XANTENNA__06923__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11549__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12407_ net1414 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
XANTENNA__07217__A1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07738__B _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13387_ net1403 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10599_ net1632 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] net837 vssd1 vssd1 vccd1
+ vccd1 _02529_ sky130_fd_sc_hd__mux2_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08965__A1 net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_105_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15126_ net1507 vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
X_12338_ net1410 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06976__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11975__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09953__B net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15057_ net1438 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
X_12269_ net1291 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__inv_2
XANTENNA__08717__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14008_ clknet_leaf_11_wb_clk_i _01772_ _00373_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06830_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] vssd1 vssd1 vccd1 vccd1
+ _02773_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13491__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ net1215 _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09480_ _02953_ net576 _05421_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08431_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XANTENNA__12029__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11215__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\] net1068
+ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ _04223_ _04234_ net847 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_4
XANTENNA__11252__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ net747 _03183_ _03184_ net1140 vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11004__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\]
+ net754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\] net1116
+ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12046__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_A _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1045_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08956__A1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__B1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1212_A team_03_WB.instance_to_wrap.core.decoder.inst\[16\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout301 _06442_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
Xfanout312 _05845_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
XANTENNA__07664__A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout334 net335 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout672_A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _06806_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
Xfanout356 _06804_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_4
XANTENNA__11186__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout367 net368 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_8
X_09816_ _05614_ _05615_ _02954_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout378 _06813_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_4
XANTENNA__10090__A _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout389 net391 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09747_ _05613_ _05688_ net576 vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06959_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\] net1146
+ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout937_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09678_ _04834_ _05577_ _05617_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09684__A2 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08629_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[102\] net940
+ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__a221o_1
XANTENNA__07695__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14782__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07790__S1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11640_ _06714_ net388 net355 net2564 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07447__A1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ net2099 net488 _06798_ net511 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13310_ net1292 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
X_10522_ net144 net1030 net1021 net1953 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07542__S1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08434__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14290_ clknet_leaf_104_wb_clk_i _02054_ _00655_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14012__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ _06037_ _06053_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13241_ net1357 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A3 _06656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input66_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ net1324 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
X_10384_ _06086_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11795__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13576__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ net1734 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14162__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07574__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12054_ _06621_ net2869 net361 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__mux2_1
XANTENNA__11703__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ net1040 net833 _06438_ net668 vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07383__B1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout890 net892 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07922__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__A1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10809__A2 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ net1341 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XANTENNA__09675__A2 _04119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ net642 _06716_ net482 net379 net2079 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a32o_1
XANTENNA__11482__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ net1416 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14626_ clknet_leaf_128_wb_clk_i _02390_ _00991_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\]
+ sky130_fd_sc_hd__dfstp_1
X_11838_ _06676_ net475 net329 net2211 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10159__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07438__A1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14557_ clknet_leaf_60_wb_clk_i _02321_ _00922_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11769_ _06602_ net479 net338 net2475 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XANTENNA__12655__A net1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13508_ net1326 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14488_ clknet_leaf_10_wb_clk_i _02252_ _00853_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[842\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10993__B2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13439_ net1424 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08399__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08938__A1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11942__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15109_ net1490 vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_2
XANTENNA__07071__C1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07610__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ net848 _04908_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__o21a_4
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07931_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\]
+ net893 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15079__1460 vssd1 vssd1 vccd1 vccd1 _15079__1460/HI net1460 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07862_ _03802_ _03803_ net811 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21o_1
XANTENNA__08571__C1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _05174_ _05338_ _05171_ _05172_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ net1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\]
+ net793 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\] net747
+ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a221o_1
XANTENNA__09115__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15206__A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09532_ _03566_ _04354_ net663 _05473_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07126__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09204__A net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _05088_ _05097_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[58\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[26\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09394_ _04415_ _05173_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_50 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08345_ net857 _04283_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21a_1
XANTENNA__08626__B1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09858__B _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout420_A _06635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1162_A net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout518_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08276_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[343\]
+ net969 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__o221a_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07227_ net720 _03152_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__o21a_4
XFILLER_0_15_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1427_A net1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07158_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[256\] net778
+ _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09051__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10736__A1 _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[577\]
+ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09085__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1107 _02786_ vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__buf_4
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
Xfanout1129 _02785_ vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_111_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11347__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09106__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ net1256 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
X_13790_ clknet_leaf_78_wb_clk_i _01554_ _00155_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07117__B1 _03043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08314__C1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12741_ net1277 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XANTENNA__07668__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12672_ net1379 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14411_ clknet_leaf_36_wb_clk_i _02175_ _00776_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08880__A3 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11623_ _06697_ net385 net353 net2510 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XANTENNA__08617__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14342_ clknet_leaf_79_wb_clk_i _02106_ _00707_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08164__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ net655 _06664_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ net114 net1028 net903 net2080 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14273_ clknet_leaf_0_wb_clk_i _02037_ _00638_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[627\]
+ sky130_fd_sc_hd__dfrtp_1
X_11485_ net2535 net399 _06776_ net511 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13224_ net1342 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
X_10436_ net305 net304 _06060_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11924__A0 _06622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ net1263 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
X_10367_ _05981_ _06089_ _06094_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12106_ net1135 net1137 _06293_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__and3_1
X_10298_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] team_03_WB.instance_to_wrap.core.pc.current_pc\[11\]
+ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and3_1
X_13086_ net1413 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12037_ net635 _06606_ net473 net368 net2293 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11257__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07356__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11554__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08339__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13988_ clknet_leaf_19_wb_clk_i _01752_ _00353_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07108__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__C1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11273__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07659__A1 team_03_WB.instance_to_wrap.core.decoder.inst\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07470__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net1271 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XANTENNA__10112__C1 _03065_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09959__A _03600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14609_ clknet_leaf_94_wb_clk_i _02373_ _00974_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08608__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12385__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ _03604_ _03728_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10966__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08061_ net1084 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\]
+ net890 _04002_ net1144 vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o311a_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07292__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07831__B2 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ net585 _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__and2_4
XFILLER_0_70_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09033__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10194__A2 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__B net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[393\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[297\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\]
+ net984 net1075 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__mux4_1
XANTENNA__08103__A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1007\]
+ net881 _03855_ net1127 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07347__B1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ net917 _04835_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__nand2_1
XANTENNA__09887__A2 _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07845_ _03779_ _03780_ _03785_ _03786_ net1107 net1130 vssd1 vssd1 vccd1 vccd1 _03787_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout370_A _06815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11464__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07661__B _03601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\]
+ net888 net1118 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__a211o_1
X_09515_ _05325_ _05327_ _05430_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08847__B1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10654__A0 net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_A net1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09446_ _05346_ _05347_ _05386_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout802_A _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _04445_ _05317_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__nor2_1
XANTENNA__11403__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11749__A3 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XANTENNA__08075__B2 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14820__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[882\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[850\]
+ net946 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09024__B1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ net499 net627 _06702_ net414 net2062 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a32o_1
XANTENNA__11906__B1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09575__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10221_ _06017_ _06021_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11382__A1 net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _03985_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__or2_1
XANTENNA__07050__A2 _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14960_ clknet_leaf_61_wb_clk_i _02712_ _01325_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__dfrtp_1
X_10083_ _02954_ _05107_ _05141_ _05082_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07338__A0 _03277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_03_WB.instance_to_wrap.core.register_file.registers_state\[937\] vssd1
+ vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ clknet_leaf_86_wb_clk_i _01675_ _00276_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[265\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07889__A1 net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14891_ clknet_leaf_44_wb_clk_i _02654_ _01256_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14200__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13842_ clknet_leaf_100_wb_clk_i _01606_ _00207_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07063__S net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__B net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13773_ clknet_leaf_104_wb_clk_i _01537_ _00138_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11437__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ _06462_ net700 vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__nor2_1
XANTENNA__11524__D net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__A0 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07105__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ net1304 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XANTENNA__14350__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ net1358 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11313__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11606_ net267 net2746 net454 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ net1249 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14325_ clknet_leaf_90_wb_clk_i _02089_ _00690_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[679\]
+ sky130_fd_sc_hd__dfrtp_1
X_11537_ net2194 net486 _06786_ net499 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XANTENNA__07813__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold409 team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\] vssd1
+ vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14256_ clknet_leaf_81_wb_clk_i _02020_ _00621_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[610\]
+ sky130_fd_sc_hd__dfrtp_1
X_11468_ net654 _06593_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__nor2_1
XANTENNA__08622__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13207_ net1418 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09566__A1 _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__S0 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _06240_ _06241_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\] net678
+ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_106_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14187_ clknet_leaf_37_wb_clk_i _01951_ _00552_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[541\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ net281 net2789 net403 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08774__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ net1420 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
XANTENNA__11983__S net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ net1318 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1109 team_03_WB.instance_to_wrap.core.register_file.registers_state\[219\] vssd1
+ vssd1 vccd1 vccd1 net2693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11125__B2 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07630_ net725 _03568_ _03569_ _03570_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a32o_1
XANTENNA__10884__B1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A2 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\]
+ net784 net1126 vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09300_ net529 _05144_ net607 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10636__A0 team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07492_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[935\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[903\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[807\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[775\]
+ net775 net1124 vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07501__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _03314_ _05161_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11223__S net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13004__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09162_ net550 _04417_ _05103_ net561 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a211o_1
XFILLER_0_28_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08113_ net1086 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\]
+ net892 net1119 vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07804__A1 net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[813\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[781\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__C _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net610 _03985_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nor2_1
XANTENNA__08532__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06841__A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold910 team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\] vssd1
+ vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 team_03_WB.instance_to_wrap.core.register_file.registers_state\[348\] vssd1
+ vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09557__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold932 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\] vssd1
+ vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold943 team_03_WB.instance_to_wrap.core.register_file.registers_state\[78\] vssd1
+ vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold954 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\] vssd1
+ vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12054__S net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11364__A1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1125_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07568__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\] vssd1
+ vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__C1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 team_03_WB.instance_to_wrap.core.register_file.registers_state\[66\] vssd1
+ vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\] vssd1
+ vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11178__B _06517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\] vssd1
+ vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _05880_ net1773 net291 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10082__B _05784_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\] net998 net938
+ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ net560 _04770_ _04817_ net665 vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11194__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[330\]
+ net1142 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21o_1
XANTENNA__10875__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07759_ net813 _03692_ net721 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12092__A2 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _02809_ vssd1 vssd1 vccd1
+ vccd1 _06380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ net584 _04830_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12440_ net1368 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08008__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15058__1439 vssd1 vssd1 vccd1 vccd1 _15058__1439/HI net1439 sky130_fd_sc_hd__conb_1
XANTENNA__11052__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12371_ net1259 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ clknet_leaf_49_wb_clk_i _01874_ _00475_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07847__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _06628_ net2629 net411 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
X_15090_ net1471 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_107_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11369__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ clknet_leaf_112_wb_clk_i _01805_ _00406_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[395\]
+ sky130_fd_sc_hd__dfrtp_1
X_11253_ net301 net711 net823 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07559__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _04739_ _05950_ _06045_ _02994_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__a211oi_1
XANTENNA__11088__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08220__A1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ net654 net707 _06527_ net697 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08678__A _04619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08508__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ team_03_WB.instance_to_wrap.core.decoder.inst\[31\] team_03_WB.instance_to_wrap.core.decoder.inst\[30\]
+ _02872_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or4_1
X_14943_ clknet_leaf_126_wb_clk_i _02698_ _01308_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11308__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ clknet_leaf_50_wb_clk_i _02637_ _01239_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07731__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ clknet_leaf_2_wb_clk_i _01589_ _00190_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[179\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13756_ clknet_leaf_119_wb_clk_i _01520_ _00121_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_10968_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[1\] net309 net684 vssd1
+ vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12083__A2 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07263__A1_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12707_ net1296 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XANTENNA__09302__A _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07495__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11830__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ clknet_leaf_87_wb_clk_i _01451_ _00052_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10899_ net271 net2085 net521 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13890__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ net1385 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09787__A1 _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11978__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12569_ net1356 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14308_ clknet_leaf_12_wb_clk_i _02072_ _00673_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold206 _02616_ vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08352__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 team_03_WB.instance_to_wrap.core.register_file.registers_state\[61\] vssd1
+ vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[48\] vssd1
+ vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11279__A net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 team_03_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1 net1823
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14239_ clknet_leaf_117_wb_clk_i _02003_ _00604_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[593\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11346__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08747__C1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08211__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08211__B2 net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 _06461_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
Xfanout719 _02864_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13494__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08800_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\] net1002
+ net923 _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__B _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09780_ _04649_ _04895_ _04956_ _05071_ net569 net563 vssd1 vssd1 vccd1 vccd1 _05722_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06992_ _02829_ _02836_ _02928_ net683 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__or4bb_2
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[964\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\] net1061
+ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11218__S net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__A1 _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_4
XANTENNA__09711__B2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[423\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[391\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[295\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[263\]
+ net980 net1074 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux4_1
XANTENNA__07846__A1_N net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07613_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\]
+ net783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\] net1158
+ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__o221a_1
X_08593_ _04478_ _04534_ net559 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_1
XANTENNA__10872__A3 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07544_ _03481_ _03485_ _03484_ net1114 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12074__A2 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11461__B _06586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11282__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[853\]
+ net762 team_03_WB.instance_to_wrap.core.register_file.registers_state\[885\] net1119
+ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o221a_1
XANTENNA__12049__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout333_A net335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ _02937_ _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09145_ net437 net430 _04323_ net550 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout500_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__D_N net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1242_A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08986__C1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09076_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[77\]
+ net962 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\] net918
+ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08027_ net1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[241\]
+ net887 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__or3_1
XANTENNA__07386__B net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 team_03_WB.instance_to_wrap.core.register_file.registers_state\[621\] vssd1
+ vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold751 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\] vssd1
+ vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _02628_ vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold773 team_03_WB.instance_to_wrap.core.register_file.registers_state\[469\] vssd1
+ vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09882__A _05596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[547\] vssd1
+ vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\] vssd1
+ vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11339__D net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ _03023_ net2539 net295 vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__mux2_1
XANTENNA__10560__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ _04867_ _04870_ net865 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_137_1629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09702__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _06633_ net2666 net375 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__mux2_1
XANTENNA__09702__B2 _04777_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__C net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ net268 net2219 net382 vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__mux2_1
X_13610_ net1297 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
X_10822_ net278 net2650 net524 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14590_ clknet_leaf_57_wb_clk_i _02354_ _00955_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_79_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08437__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13541_ net1329 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08364__S1 net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11371__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10753_ net324 net602 vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11812__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13472_ net1327 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XANTENNA_input96_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ _05429_ _06313_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15211_ net1577 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XANTENNA__11798__S net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13579__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ net1389 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15142_ net1523 vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ net1364 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _06615_ net2677 net409 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XANTENNA__11099__A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15073_ net1454 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
X_12285_ net1382 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ clknet_leaf_35_wb_clk_i _01788_ _00389_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[378\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ net506 net631 _06685_ net416 net2715 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net694 net709 net298 vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__or3b_1
XFILLER_0_101_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10551__A2 _06293_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10118_ _05960_ net2872 _05947_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ _06625_ net2555 net424 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11265__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14926_ clknet_leaf_123_wb_clk_i _02681_ _01291_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_10049_ net7 net1036 net908 net2876 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08901__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14857_ clknet_leaf_42_wb_clk_i net1851 _01222_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10877__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_114_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13808_ clknet_leaf_83_wb_clk_i _01572_ _00173_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14788_ clknet_leaf_56_wb_clk_i _02552_ _01153_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11264__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13739_ clknet_leaf_27_wb_clk_i _01503_ _00104_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07468__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09967__A _03788_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ net1124 _03198_ _03199_ net1110 vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11016__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13489__A net1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[883\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[851\]
+ net754 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11501__S net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07487__A _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08968__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08432__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08983__A2 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _05834_ _05841_ _05833_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10790__A2 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_888 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11159__D net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout505 _06448_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout516 net520 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_2
X_09832_ net580 _04711_ _04821_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__o31a_1
Xfanout538 _06298_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XANTENNA__08291__S0 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 _03106_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07943__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ net358 _05463_ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08111__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[517\] net790
+ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout283_A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[196\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[228\] net923
+ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057__1438 vssd1 vssd1 vccd1 vccd1 _15057__1438/HI net1438 sky130_fd_sc_hd__conb_1
X_09694_ _05196_ _05203_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09160__A2 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07950__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\]
+ net1003 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\] net939
+ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout450_A _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__A1 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _04512_ _04517_ net868 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07527_ _03467_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__B1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07458_ net739 _03398_ _03399_ net801 vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a31o_1
XANTENNA__08671__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08671__B2 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07389_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\] net768
+ _02871_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11411__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14561__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ net440 net432 _05068_ net546 vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__o31a_1
XFILLER_0_66_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09059_ _04999_ _05000_ net1062 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08005__B _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ _06546_ net2560 net364 vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__mux2_1
Xhold570 team_03_WB.instance_to_wrap.core.register_file.registers_state\[827\] vssd1
+ vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 team_03_WB.instance_to_wrap.core.register_file.registers_state\[439\] vssd1
+ vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold592 team_03_WB.instance_to_wrap.core.register_file.registers_state\[364\] vssd1
+ vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ net2283 net427 _06584_ net500 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10533__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A1 _06499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09117__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ net1299 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1270 team_03_WB.instance_to_wrap.core.register_file.registers_state\[210\] vssd1
+ vssd1 vccd1 vccd1 net2854 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09551__S net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1281 team_03_WB.instance_to_wrap.ADR_I\[30\] vssd1 vssd1 vccd1 vccd1 net2865
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ _06479_ net2521 net374 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__mux2_1
X_14711_ clknet_leaf_11_wb_clk_i _02475_ _01076_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1292 team_03_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1 net2876
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ clknet_leaf_100_wb_clk_i _02406_ _01007_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[996\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _06453_ net2178 net381 vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11246__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__S1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ _06410_ _06411_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__a21oi_4
X_14573_ clknet_leaf_106_wb_clk_i _02337_ _00938_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[927\]
+ sky130_fd_sc_hd__dfrtp_1
X_11785_ net2608 _06618_ net335 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__mux2_1
XANTENNA__11532__D net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13659__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11797__A1 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ net1273 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10736_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] _05659_ net603 vssd1
+ vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ net1331 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _02765_ _06305_ _06306_ _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11549__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11321__S net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ net1344 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
X_13386_ net1331 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ net1646 team_03_WB.instance_to_wrap.CPU_DAT_O\[31\] net835 vssd1 vssd1 vccd1
+ vccd1 _02530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15125_ net1506 vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_2
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
X_12337_ net1303 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12941__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15056_ net1437 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_120_162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12268_ net1300 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14007_ clknet_leaf_75_wb_clk_i _01771_ _00372_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ net298 net2562 net491 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__mux2_1
XANTENNA__11557__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net1598 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10524__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__A1 _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07246__S net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11991__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14909_ clknet_leaf_39_wb_clk_i _00003_ _01274_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07689__C1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07153__A1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08430_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[666\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\] net918
+ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ net857 _04299_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11788__A1 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ net1143 _03252_ _03253_ net816 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o31a_1
XANTENNA__14584__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09697__A _03866_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _04228_ _04233_ net870 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10460__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07243_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[584\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[616\] net730
+ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o221a_1
XANTENNA__11231__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07174_ net806 _03112_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08106__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07010__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07613__C1 net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1038_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout302 _06438_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XANTENNA_fanout498_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12062__S net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10515__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1205_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__buf_4
XANTENNA__11712__A1 _06409_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__B1 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout346 net347 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__buf_6
X_09815_ _02954_ _05587_ _05749_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a211o_4
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__B _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 _06817_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_6
XANTENNA__10090__B _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout379 net380 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_6
XFILLER_0_96_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout665_A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _05084_ _05086_ _05117_ _05119_ net556 net572 vssd1 vssd1 vccd1 vccd1 _05688_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06958_ net805 _02896_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09677_ _03391_ _04119_ net664 _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07144__A1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout832_A _06386_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06889_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] _02820_ vssd1 vssd1 vccd1
+ vccd1 _02831_ sky130_fd_sc_hd__and2_1
XANTENNA__11406__S net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08628_ _04568_ _04569_ net852 vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o21a_1
XANTENNA__13801__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14927__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11228__A0 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ net1055 _04497_ _04500_ net863 vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11570_ net637 net706 net267 net697 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__and4_1
XANTENNA__08644__A1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10521_ net145 net1024 net1022 net1783 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07852__C1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13240_ net1369 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
X_10452_ net305 net304 _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__and3_1
XANTENNA__08016__A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11400__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13171_ net1264 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
X_10383_ _05994_ _06085_ _05996_ _05992_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12761__A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06958__A1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12122_ net1668 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07080__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input59_A gpio_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ _06469_ net2870 net361 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__mux2_1
XANTENNA__10506__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ net2423 net427 _06574_ net515 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a22o_1
XANTENNA__07293__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07383__A1 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__C1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__B1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net882 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13592__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout891 net892 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_2
XANTENNA__07590__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ net1344 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11316__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A3 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ net637 _06715_ net478 net379 net2171 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12886_ net1344 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11219__A0 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ net654 _06675_ net475 net329 net1738 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a32o_1
X_14625_ clknet_leaf_134_wb_clk_i _02389_ _00990_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[979\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08096__C1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14556_ clknet_leaf_127_wb_clk_i _02320_ _00921_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11768_ _06601_ net482 net338 net2446 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10442__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09310__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ net1324 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
X_10719_ _05596_ net601 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ clknet_leaf_75_wb_clk_i _02251_ _00852_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\]
+ sky130_fd_sc_hd__dfrtp_1
X_11699_ _06741_ net390 net347 net2170 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10993__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13438_ net1314 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15056__1437 vssd1 vssd1 vccd1 vccd1 _15056__1437/HI net1437 sky130_fd_sc_hd__conb_1
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08399__B1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13369_ net1326 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XANTENNA__09060__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09060__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06949__A1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A1 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07071__B1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15108_ net1489 vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_2
XANTENNA__11287__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15039_ clknet_leaf_33_wb_clk_i _02759_ _01404_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__dfrtp_1
X_07930_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\]
+ net768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\] net729
+ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07861_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[667\]
+ net729 _03791_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ _05541_ _05500_ _05518_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3b_1
XANTENNA__08571__B1 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[683\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[651\]
+ net771 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__mux2_1
XANTENNA__08596__A _02954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09531_ _03566_ _04354_ net541 vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09746__S0 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07931__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11226__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10130__A0 _04415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _05397_ _05403_ net581 vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08413_ net440 net432 _04354_ net551 vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _05318_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or3b_2
XFILLER_0_87_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_62 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ net851 _04284_ _04285_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07429__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06844__A net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__C _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12057__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ net854 _04215_ _04216_ _04214_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout413_A net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07226_ net1138 _03159_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09051__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07157_ net1189 team_03_WB.instance_to_wrap.core.register_file.registers_state\[288\]
+ net879 _02872_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12581__A net1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1322_A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07088_ net746 _03028_ _03029_ net1156 vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout782_A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1119 net1120 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_4
XANTENNA__11697__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ _04150_ _04269_ _04326_ _04386_ net568 net564 vssd1 vssd1 vccd1 vccd1 _05671_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07117__A1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12740_ net1306 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08865__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12671_ net1374 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14410_ clknet_leaf_3_wb_clk_i _02174_ _00775_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[764\]
+ sky130_fd_sc_hd__dfrtp_1
X_11622_ _06696_ net385 net353 net2609 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XANTENNA__08617__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14341_ clknet_leaf_107_wb_clk_i _02105_ _00706_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[695\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11621__B1 net356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ net2360 net487 _06791_ net501 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ net125 net1028 net903 net1717 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14272_ clknet_leaf_133_wb_clk_i _02036_ _00637_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[626\]
+ sky130_fd_sc_hd__dfrtp_1
X_11484_ net637 net706 _06550_ net824 vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ net1403 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
Xwire588 _04861_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_4
XFILLER_0_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ _06253_ _06254_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] net679
+ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09042__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10727__A2 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07585__A team_03_WB.instance_to_wrap.core.decoder.inst\[24\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ net1346 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08180__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10366_ _05981_ _06089_ _06094_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ _06799_ net482 net446 net2371 vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13085_ net1381 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
X_10297_ team_03_WB.instance_to_wrap.core.pc.current_pc\[10\] _06138_ vssd1 vssd1
+ vccd1 vccd1 _06139_ sky130_fd_sc_hd__and2_1
X_12036_ _06775_ net478 net367 net2476 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a22o_1
XANTENNA__11688__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06929__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07524__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09305__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ clknet_leaf_24_wb_clk_i _01751_ _00352_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[341\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11273__C net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ net1258 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
XANTENNA__07659__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11860__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09959__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12869_ net1274 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11570__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08608__A1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ clknet_leaf_80_wb_clk_i _02372_ _00973_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__08355__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09040__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11612__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14539_ clknet_leaf_37_wb_clk_i _02303_ _00904_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08084__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10966__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08060_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\]
+ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__or2_1
XANTENNA__07292__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07011_ net529 _02944_ _02948_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__and4_2
XANTENNA__13497__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09033__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10914__A _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__D_N net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07926__C net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_942 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[489\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__o221a_1
XANTENNA__11448__C net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07913_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\]
+ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__and2_1
XANTENNA__11679__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ _02795_ _02796_ net958 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07347__A1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07844_ _03781_ _03782_ net738 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__mux2_1
XANTENNA__06839__A team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07775_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\]
+ net874 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout363_A net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _05327_ _05430_ _05325_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__o21a_1
XANTENNA__08847__A1 net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ _05346_ _05347_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11851__A0 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout530_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_A net1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _04445_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__and2_1
XANTENNA__08265__S net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10808__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11603__A0 _06536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ net550 _04237_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07807__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10096__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10957__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08258_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\]
+ net948 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08480__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout997_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07209_ net1151 _03149_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09024__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08189_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[435\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[403\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[307\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[275\]
+ net950 net1065 vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09096__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07609__S net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ _06057_ _06059_ _06022_ _06024_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a211o_1
XANTENNA__07035__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _04178_ team_03_WB.instance_to_wrap.core.pc.current_pc\[17\] net674 vssd1
+ vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _05768_ _05784_ _05798_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__and3_1
X_13910_ clknet_leaf_84_wb_clk_i _01674_ _00275_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[264\]
+ sky130_fd_sc_hd__dfrtp_1
X_14890_ clknet_leaf_43_wb_clk_i _02653_ _01255_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13841_ clknet_leaf_96_wb_clk_i _01605_ _00206_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[195\]
+ sky130_fd_sc_hd__dfrtp_1
X_15055__1436 vssd1 vssd1 vccd1 vccd1 _15055__1436/HI net1436 sky130_fd_sc_hd__conb_1
XFILLER_0_74_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12095__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ clknet_leaf_7_wb_clk_i _01536_ _00137_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10984_ net1245 net828 vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__or2_4
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08964__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ net1259 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__S0 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ net1340 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11605_ _06545_ net2518 net454 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12585_ net1248 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ net628 _06646_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__and2_1
X_14324_ clknet_leaf_92_wb_clk_i _02088_ _00689_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ clknet_leaf_98_wb_clk_i _02019_ _00620_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ net2410 net397 _06769_ net501 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
X_13206_ net1338 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
X_10418_ net285 _06140_ _06238_ net678 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o31a_1
XANTENNA__09110__S1 net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14186_ clknet_leaf_2_wb_clk_i _01950_ _00551_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[540\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08204__A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ _06449_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__or2_4
XANTENNA__07577__A1 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08774__B1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ net1314 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_10349_ _02771_ _06148_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13068_ net1305 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
XANTENNA__11125__A2 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ net616 _06580_ net458 net365 net2461 vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07560_ net1187 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\] team_03_WB.instance_to_wrap.core.decoder.inst\[22\]
+ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__o221a_1
XANTENNA__12086__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11428__A3 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10636__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11833__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07491_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11504__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ _04532_ _05169_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09161_ net437 net429 _04532_ net544 vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__o31a_1
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[698\]
+ net875 vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09092_ net1199 _05030_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08813__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ net1203 _02821_ _03107_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09006__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\] vssd1
+ vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09006__B2 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold911 team_03_WB.instance_to_wrap.core.register_file.registers_state\[120\] vssd1
+ vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold922 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\] vssd1
+ vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12010__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08214__C1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\] vssd1
+ vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold944 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\] vssd1
+ vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold955 net202 vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11364__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__B1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\] vssd1
+ vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 team_03_WB.instance_to_wrap.core.register_file.registers_state\[857\] vssd1
+ vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09994_ _05879_ net2249 net287 vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1020_A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\] vssd1
+ vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11178__C _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[325\] vssd1
+ vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1118_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10082__C _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\]
+ net974 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout480_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A _02993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14518__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _02831_ _02929_ _02935_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__or3b_4
XFILLER_0_97_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11194__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ net1166 team_03_WB.instance_to_wrap.core.register_file.registers_state\[362\]
+ net872 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__and3_1
XANTENNA__10875__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout745_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07758_ net813 _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12077__B1 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10088__C1 _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10627__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11824__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09428_ _04832_ _05368_ _05369_ _05364_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09359_ _05291_ _05296_ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__or3_1
XFILLER_0_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08048__A2 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13692__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ net1412 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08453__C1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07351__S0 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ _06627_ net2816 net410 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__mux2_1
XANTENNA__07847__B net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12001__A0 _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14040_ clknet_leaf_118_wb_clk_i _01804_ _00405_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09548__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ net507 net630 _06693_ net416 net2531 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a32o_1
XANTENNA__11369__B _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14048__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__A1 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10203_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] _05950_ vssd1 vssd1 vccd1
+ vccd1 _06045_ sky130_fd_sc_hd__nor2_1
XANTENNA__08756__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11183_ net2188 net419 _06672_ net513 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a22o_1
XANTENNA__10563__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08959__A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _03565_ _05974_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nor2_1
XANTENNA__07863__A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A gpio_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08508__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14942_ clknet_leaf_39_wb_clk_i _02697_ _01307_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10065_ team_03_WB.instance_to_wrap.core.decoder.inst\[24\] net1139 net1178 team_03_WB.instance_to_wrap.core.decoder.inst\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14873_ clknet_leaf_50_wb_clk_i _02636_ _01238_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12068__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ clknet_leaf_132_wb_clk_i _01588_ _00189_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10618__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__B1 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ clknet_leaf_28_wb_clk_i _01519_ _00120_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[109\]
+ sky130_fd_sc_hd__dfrtp_1
X_10967_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[1\] net306 vssd1 vssd1
+ vccd1 vccd1 _06547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11324__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ net1364 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XANTENNA__07495__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08692__C1 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10898_ _06488_ _06489_ _06490_ net586 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__o211a_1
X_13686_ clknet_leaf_84_wb_clk_i _01450_ _00051_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07103__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ net1375 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA__08039__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09787__A2 _05508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ net1370 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XANTENNA__08995__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14307_ clknet_leaf_18_wb_clk_i _02071_ _00672_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11519_ _06632_ net2501 net395 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ net1259 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold207 team_03_WB.instance_to_wrap.core.register_file.registers_state\[28\] vssd1
+ vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_03_WB.instance_to_wrap.ADR_I\[17\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 net234 vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ clknet_leaf_49_wb_clk_i _02002_ _00603_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[592\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11279__B _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11346__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11994__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ clknet_leaf_112_wb_clk_i _01933_ _00534_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07014__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10554__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__A _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ net1016 net821 _02825_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__nor4b_1
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[804\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\]
+ net975 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1280 net1295 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_4
XANTENNA__09711__A2 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08661_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[455\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\] net1074
+ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a221o_1
Xfanout1291 net1295 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_4
X_07612_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[793\] net798
+ _03548_ net1113 vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08592_ _04505_ _04533_ net551 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ net1124 _03483_ net1160 vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07370__A1_N net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09475__A1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07486__A0 _03425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11282__A1 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07474_ _03411_ _03415_ net1138 vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11821__A3 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__A_N _05654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ _03429_ _04032_ net438 _05146_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__or4_2
XANTENNA__07013__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1068_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ net546 _04179_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07948__A net1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11034__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08770__C _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08986__B1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ net933 _05015_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12065__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1235_A net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15054__1435 vssd1 vssd1 vccd1 vccd1 _15054__1435/HI net1435 sky130_fd_sc_hd__conb_1
X_08026_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[81\]
+ net760 team_03_WB.instance_to_wrap.core.register_file.registers_state\[113\] net728
+ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold730 team_03_WB.instance_to_wrap.core.register_file.registers_state\[110\] vssd1
+ vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[11\] vssd1 vssd1 vccd1
+ vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout695_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[736\] vssd1
+ vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\] vssd1
+ vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\] vssd1
+ vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1402_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 team_03_WB.instance_to_wrap.core.register_file.registers_state\[506\] vssd1
+ vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\] vssd1
+ vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07683__A net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09977_ net590 net1870 net294 vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout862_A _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07961__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11409__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net860 _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08859_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[928\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[800\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[768\]
+ net986 net1074 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_58_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ _06536_ net2395 net382 vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10821_ _06423_ _06425_ net587 vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__o21a_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ net1326 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
X_10752_ team_03_WB.instance_to_wrap.core.pc.current_pc\[6\] net602 vssd1 vssd1 vccd1
+ vccd1 _06369_ sky130_fd_sc_hd__or2_1
XANTENNA__07477__B1 net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11371__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ net1393 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10683_ _06321_ net525 _06324_ net530 net2810 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a32o_1
XFILLER_0_82_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ net911 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__clkbuf_1
X_12422_ net1412 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input89_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15141_ net1522 vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
XFILLER_0_51_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ net1290 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ _06614_ net2753 net411 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__mux2_1
X_15072_ net1453 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_121_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11099__B net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ net1350 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14023_ clknet_leaf_66_wb_clk_i _01787_ _00388_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\]
+ sky130_fd_sc_hd__dfrtp_1
X_11235_ _06405_ net716 net826 vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__and3_1
XANTENNA__10536__B1 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11879__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ net2234 net418 _06661_ net503 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11319__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10117_ _05954_ _05955_ _03065_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11097_ net828 net299 vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10839__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[22\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ net8 net1034 _05907_ net1823 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__o22a_1
X_14925_ clknet_leaf_124_wb_clk_i _02680_ _01290_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__A1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12939__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1002\] vssd1
+ vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08901__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14856_ clknet_leaf_42_wb_clk_i net1803 _01221_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09313__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13807_ clknet_leaf_99_wb_clk_i _01571_ _00172_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[161\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14787_ clknet_leaf_55_wb_clk_i _02551_ _01152_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11999_ _06523_ net2331 net451 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07468__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ clknet_leaf_4_wb_clk_i _01502_ _00103_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11281__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13669_ clknet_leaf_106_wb_clk_i _01433_ _00034_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11016__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[787\]
+ net754 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08968__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__B _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14363__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _05834_ _05841_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and2_2
XFILLER_0_50_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10527__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout517 net520 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
X_09831_ net579 _04711_ net665 _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a22o_1
Xfanout528 _06322_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_2
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07943__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08291__S1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11229__S net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ _04327_ _05073_ _05702_ _05703_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__a211o_1
X_06974_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[645\]
+ net770 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\] net743
+ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__o221a_1
X_08713_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[68\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[100\] net939
+ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a221o_1
X_09693_ _05276_ _05279_ _05198_ _05207_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_59_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ net922 _04584_ _04585_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06847__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09223__A _04503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ net1211 _04515_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_1696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_A _04075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07526_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[710\]
+ net795 team_03_WB.instance_to_wrap.core.register_file.registers_state\[742\] net731
+ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07457_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\]
+ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12584__A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1352_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout708_A _06461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11007__B2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14706__CLK clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07388_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[287\] net791
+ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11558__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__inv_2
XANTENNA__09081__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[623\] net942
+ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08009_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[849\]
+ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_664 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold560 net225 vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 team_03_WB.instance_to_wrap.core.register_file.registers_state\[55\] vssd1
+ vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08187__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\] vssd1
+ vssd1 vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net627 _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__nor2_1
Xhold593 team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\] vssd1
+ vssd1 vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08302__A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06867__C_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09687__A1 _04829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ net1272 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XANTENNA__07147__C1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1260 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[9\] vssd1 vssd1 vccd1
+ vccd1 net2844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1271 team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\] vssd1
+ vssd1 vccd1 vccd1 net2855 sky130_fd_sc_hd__dlygate4sd3_1
X_14710_ clknet_leaf_116_wb_clk_i _02474_ _01075_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.decoder.inst\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11922_ _06621_ net2854 net373 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__mux2_1
Xhold1282 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\] vssd1
+ vssd1 vccd1 vccd1 net2866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] vssd1 vssd1 vccd1 vccd1
+ net2877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08895__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14236__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__A _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ clknet_leaf_102_wb_clk_i _02405_ _01006_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[995\]
+ sky130_fd_sc_hd__dfstp_1
X_11853_ _06446_ net2216 net384 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10049__A2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__A1 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ net689 _05563_ _06401_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ net2319 _06617_ net334 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__mux2_1
X_14572_ clknet_leaf_7_wb_clk_i _02336_ _00937_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\]
+ sky130_fd_sc_hd__dfrtp_1
X_15169__1550 vssd1 vssd1 vccd1 vccd1 _15169__1550/HI net1550 sky130_fd_sc_hd__conb_1
XFILLER_0_68_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13523_ net1278 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
X_10735_ net2089 net530 net525 _06359_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11602__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13454_ net1393 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
X_10666_ net1137 _06307_ _06302_ team_03_WB.instance_to_wrap.core.ru.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07870__B1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10206__C1 _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11549__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06923__C net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ net1264 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
X_13385_ net1309 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_10597_ net1134 team_03_WB.instance_to_wrap.core.d_hit team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ _06281_ net838 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ net1505 vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_2
XFILLER_0_51_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
X_12336_ net1428 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06976__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12267_ net1253 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__inv_2
X_15055_ net1436 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__10509__B1 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11218_ net299 net2778 net491 vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__mux2_1
X_14006_ clknet_leaf_86_wb_clk_i _01770_ _00371_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09308__A _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ net1587 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07925__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ net495 net647 _06651_ net417 net1925 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a32o_1
XANTENNA__15011__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09678__A1 _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08866__B _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14908_ clknet_leaf_38_wb_clk_i _00002_ _01273_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07689__B1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11485__B2 net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__A1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14839_ clknet_leaf_57_wb_clk_i _02603_ _01204_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_1
X_15053__1434 vssd1 vssd1 vccd1 vccd1 _15053__1434/HI net1434 sky130_fd_sc_hd__conb_1
XANTENNA__10189__A _03460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12029__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ net851 _04300_ _04301_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__or3_1
XANTENNA__08638__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08882__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ net1176 team_03_WB.instance_to_wrap.core.register_file.registers_state\[861\]
+ net765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\] net1154
+ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08291_ _04229_ _04230_ _04231_ _04232_ net856 net932 vssd1 vssd1 vccd1 vccd1 _04233_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09697__B _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07310__C1 net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11512__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ net1184 team_03_WB.instance_to_wrap.core.register_file.registers_state\[712\]
+ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__or2_1
XANTENNA__10460__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13753__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ net801 _03113_ _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07613__B1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07010__B net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout303 _06422_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_2
XANTENNA__09218__A _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout314 _05388_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_4
Xfanout325 _05355_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07664__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_A net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _06810_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09814_ _05754_ _05755_ _05752_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__or3b_1
Xfanout347 _06806_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11186__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 _04831_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__clkbuf_4
Xfanout369 net370 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1100_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__C _05659_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _05213_ _05235_ _05275_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__nand3_1
XANTENNA__09669__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout560_A _03064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ net808 _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__and3_1
XANTENNA__12579__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_A _06457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ _03391_ _04119_ net542 vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o21ai_1
X_06888_ _02822_ _02823_ _02827_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__or4_1
XANTENNA__11476__B2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08341__A1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ net1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[134\]
+ net979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[166\] net940
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_A net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08629__C1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08558_ _04498_ _04499_ net1208 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07509_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\] net1148
+ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_135_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08489_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[59\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[27\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09841__A1 _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11422__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ net146 net1023 net1019 net2005 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13203__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__B _04475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07852__B1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10451_ _06135_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13170_ net1422 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
XANTENNA__07604__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10382_ team_03_WB.instance_to_wrap.core.pc.current_pc\[18\] _06144_ vssd1 vssd1
+ vccd1 vccd1 _06211_ sky130_fd_sc_hd__xor2_1
XANTENNA__08801__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12121_ net1709 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07080__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15034__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _06454_ net2761 net361 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__mux2_1
Xhold390 team_03_WB.instance_to_wrap.CPU_DAT_I\[15\] vssd1 vssd1 vccd1 vccd1 net1974
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11377__B net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07368__C1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ net275 net658 net705 net826 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__and4_1
XANTENNA__11703__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08580__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09109__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__clkbuf_8
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout892 net901 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11393__A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ net1368 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
XANTENNA__11467__B2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\] vssd1
+ vssd1 vccd1 vccd1 net2674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_137_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11905_ net632 _06714_ net470 net380 net2184 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a32o_1
X_12885_ net1262 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14624_ clknet_leaf_134_wb_clk_i _02388_ _00989_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11836_ net653 _06674_ net468 net329 net1936 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14555_ clknet_leaf_28_wb_clk_i _02319_ _00920_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08096__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ _06599_ net480 net338 net2359 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XANTENNA__09832__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ net1310 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XANTENNA__13113__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\] net600 vssd1 vssd1 vccd1
+ vccd1 _06350_ sky130_fd_sc_hd__or2_1
XANTENNA__10442__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14486_ clknet_leaf_85_wb_clk_i _02250_ _00851_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08207__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11698_ _06740_ net387 net344 net2383 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07111__A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13437_ net1314 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10649_ team_03_WB.instance_to_wrap.core.decoder.inst\[12\] team_03_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ net841 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
XANTENNA__08399__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__B1 _05531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ net1326 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06949__A2 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1488 vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_2
XANTENNA__07071__A1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319_ net1377 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
X_13299_ net1394 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
X_15038_ clknet_leaf_62_wb_clk_i _02758_ _01403_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11287__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__C1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07860_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\] net780
+ net748 _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08571__A1 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07791_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[555\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[523\]
+ net772 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__mux2_1
XANTENNA__12399__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09530_ net581 _05471_ net358 vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07126__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__A1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _05399_ _05402_ net573 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ net848 _04340_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__o21ba_4
X_09392_ _04382_ _05312_ _05319_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09501__A _03823_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[213\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\] net935
+ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08626__A2 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10969__B1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[215\]
+ net970 team_03_WB.instance_to_wrap.core.register_file.registers_state\[247\] net937
+ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__o221a_1
XANTENNA__07834__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07225_ net1130 _03162_ _03164_ _03166_ net720 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o41a_1
XFILLER_0_6_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1050_A _02791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A _06718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1148_A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[384\] net778
+ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11394__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07062__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07087_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[673\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__or3_1
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1315_A net1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14081__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1109 _02786_ vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07365__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[816\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[784\]
+ net784 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11417__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07770__C1 net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _04210_ _05014_ _05071_ _04895_ net559 net574 vssd1 vssd1 vccd1 vccd1 _05670_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11449__B2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__A2 _03058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _05084_ _05089_ _05091_ _05098_ net566 net562 vssd1 vssd1 vccd1 vccd1 _05601_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11941__A _02793_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12670_ net1385 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11621_ _06695_ net386 net356 net2299 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14340_ clknet_leaf_12_wb_clk_i _02104_ _00705_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ net651 _06662_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08027__A net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ net2252 net1028 net903 net2135 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14271_ clknet_leaf_121_wb_clk_i _02035_ _00636_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\]
+ sky130_fd_sc_hd__dfrtp_1
X_11483_ net515 net635 _06606_ net400 net2414 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input71_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ net1429 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
X_10434_ net284 _06138_ _06250_ net679 vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__o31a_1
XANTENNA__07866__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire589 _04679_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__buf_4
XANTENNA__14424__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10365_ team_03_WB.instance_to_wrap.core.pc.current_pc\[20\] _06145_ team_03_WB.instance_to_wrap.core.pc.current_pc\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07585__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ net1276 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12104_ _06798_ net478 net445 net2162 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a22o_1
X_13084_ net1350 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
X_10296_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] team_03_WB.instance_to_wrap.core.pc.current_pc\[8\]
+ _06136_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12035_ net636 _06604_ net475 net367 net2153 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a32o_1
XANTENNA__14574__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11327__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09728__S1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ clknet_leaf_130_wb_clk_i _01750_ _00351_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08305__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09502__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12101__A2 _06675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07106__A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10112__A1 _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12937_ net1252 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12868_ net1306 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__B net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607_ clknet_leaf_98_wb_clk_i _02371_ _00972_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08069__B1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ _06649_ net467 net328 net2362 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12799_ net1376 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14538_ clknet_leaf_3_wb_clk_i _02302_ _00903_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__S net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10966__A3 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09018__C1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07292__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14469_ clknet_leaf_122_wb_clk_i _02233_ _00834_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07010_ net1018 net583 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09569__B1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08371__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11376__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08792__A1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ net1235 team_03_WB.instance_to_wrap.core.register_file.registers_state\[329\]
+ net984 team_03_WB.instance_to_wrap.core.register_file.registers_state\[361\] net1075
+ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11448__D net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[879\]
+ net881 _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08892_ net580 net358 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148__1529 vssd1 vssd1 vccd1 vccd1 _15148__1529/HI net1529 sky130_fd_sc_hd__conb_1
X_07843_ _03783_ _03784_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13941__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07774_ net1084 net890 team_03_WB.instance_to_wrap.core.register_file.registers_state\[524\]
+ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__o21a_1
XANTENNA__09930__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09513_ _05435_ _05453_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__or2_1
XANTENNA__11300__A0 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12857__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1098_A net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _05371_ _05385_ _05370_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09231__A _03314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09375_ _05160_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12068__S net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08326_ net440 net432 _04267_ net545 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__o31a_1
XANTENNA__07807__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10096__B _05429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08257_ net929 _04197_ _04198_ net850 vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__o211a_1
XANTENNA__08480__B1 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__B _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1432_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07208_ net1106 _03147_ _03148_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08281__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[467\]
+ net947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__o221a_1
XFILLER_0_43_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout892_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07139_ _03077_ _03080_ net815 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09980__A0 _03103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _03139_ _05990_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _05918_ _05923_ _05924_ _02831_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__a211o_2
XFILLER_0_96_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13840_ clknet_leaf_82_wb_clk_i _01604_ _00205_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[194\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10893__A2 _06486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06864__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12095__A1 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ clknet_leaf_36_wb_clk_i _01535_ _00136_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08299__B1 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ net1245 net828 vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12722_ net1419 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09141__A net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06944__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ net1301 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ net268 net2686 net454 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ net1352 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07274__A1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14323_ clknet_leaf_109_wb_clk_i _02087_ _00688_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07274__B2 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ net2481 net489 _06785_ net516 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14254_ clknet_leaf_69_wb_clk_i _02018_ _00619_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[608\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11466_ net651 _06591_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11358__B1 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ net1269 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
X_10417_ _05925_ _05945_ _06067_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a211o_1
X_14185_ clknet_leaf_59_wb_clk_i _01949_ _00550_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[539\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11397_ net649 _06459_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__or2_4
XFILLER_0_104_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12007__A net1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ net1428 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10348_ _06107_ _06109_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__xor2_1
XANTENNA__10581__B2 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10750__A _05730_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _03822_ _06117_ _06114_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13067_ net1275 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
XANTENNA__08526__A1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ net621 _06579_ net461 net365 net2131 vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07762__C net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12086__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ clknet_leaf_94_wb_clk_i _01733_ _00334_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07490_ net1101 team_03_WB.instance_to_wrap.core.register_file.registers_state\[967\]
+ net797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[999\] net1126
+ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07501__A2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ net544 _04476_ _05101_ net555 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08890__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__A0 net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08111_ net1175 team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\]
+ net875 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ net933 _05032_ _05031_ net1056 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11520__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ net717 _03962_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_1299 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 team_03_WB.instance_to_wrap.core.register_file.registers_state\[155\] vssd1
+ vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold912 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\] vssd1
+ vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07017__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold923 team_03_WB.instance_to_wrap.core.register_file.registers_state\[918\] vssd1
+ vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold934 team_03_WB.instance_to_wrap.core.register_file.registers_state\[514\] vssd1
+ vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold945 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\] vssd1
+ vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09962__A0 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold956 team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\] vssd1
+ vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08765__A1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07568__A2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\] vssd1
+ vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold978 team_03_WB.instance_to_wrap.core.register_file.registers_state\[780\] vssd1
+ vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05878_ net1820 net287 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__mux2_1
Xhold989 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\] vssd1
+ vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ net1047 team_03_WB.instance_to_wrap.core.register_file.registers_state\[715\]
+ net1002 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\] net923
+ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__a221o_1
X_08875_ net559 _04770_ net542 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11875__D_N net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07826_ _03764_ _03767_ net812 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11194__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12077__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09478__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ net1153 _03697_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout640_A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout738_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07688_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\] net1115
+ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__o221a_1
XANTENNA__08150__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07180__S net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _04476_ _05081_ _05126_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__or3b_1
XFILLER_0_133_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout905_A _06285_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13837__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _05298_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11588__A0 _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08309_ net864 _04250_ _04245_ net843 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08008__C net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A2 net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ _06505_ net2722 net411 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__mux2_1
XANTENNA__07351__S1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ net1243 net833 net302 net669 vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__and4_1
XFILLER_0_107_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11369__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10012__A0 _03059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08756__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10202_ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] net672 vssd1 vssd1 vccd1
+ vccd1 _06044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ net639 _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11760__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _03565_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08508__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ clknet_leaf_126_wb_clk_i _02696_ _01306_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input34_A gpio_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ team_03_WB.instance_to_wrap.core.decoder.inst\[11\] team_03_WB.instance_to_wrap.core.decoder.inst\[10\]
+ net1240 net1245 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or4_1
XANTENNA__11512__A0 _06519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14872_ clknet_leaf_37_wb_clk_i net1728 _01237_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.wb.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A2 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09502__A2_N net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13823_ clknet_leaf_121_wb_clk_i _01587_ _00188_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14612__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11605__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10079__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__A1 net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13754_ clknet_leaf_22_wb_clk_i _01518_ _00119_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10966_ net509 net593 net263 net522 net1865 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a32o_1
XFILLER_0_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12705_ net1290 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07495__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ clknet_leaf_89_wb_clk_i _01449_ _00050_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_10897_ net685 _05821_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12636_ net1341 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XANTENNA__11579__A0 _06418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08914__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15147__1528 vssd1 vssd1 vccd1 vccd1 _15147__1528/HI net1528 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10745__A _05706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ net1413 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ clknet_leaf_127_wb_clk_i _02070_ _00671_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[660\]
+ sky130_fd_sc_hd__dfrtp_1
X_11518_ net263 net2588 net396 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__mux2_1
X_12498_ net1412 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
Xhold208 net135 vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_830 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold219 _02620_ vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14237_ clknet_leaf_68_wb_clk_i _02001_ _00602_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[591\]
+ sky130_fd_sc_hd__dfrtp_1
X_11449_ net2614 net399 _06763_ net516 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10003__A0 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11279__C net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08747__A1 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14168_ clknet_leaf_119_wb_clk_i _01932_ _00533_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[522\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__B1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07955__C1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ net1378 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ clknet_leaf_110_wb_clk_i _01863_ _00464_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06990_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__B _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__A0 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1270 net1433 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_4
Xfanout1281 net1283 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_4
X_08660_ net1051 team_03_WB.instance_to_wrap.core.register_file.registers_state\[327\]
+ net1005 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__a221o_1
XANTENNA__09711__A3 _05041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1292 net1294 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_4
X_07611_ net1113 _03551_ _03552_ net1127 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08591_ net440 net432 _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11515__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07542_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[422\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[390\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[294\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[262\]
+ net775 net1124 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux4_1
XANTENNA__11806__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07473_ _03413_ _03414_ net1153 vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11282__A2 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09212_ _03391_ _03428_ _05152_ net605 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__a31o_1
XANTENNA__10490__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07238__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ net439 net431 _04984_ net552 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__o31a_1
XANTENNA__11034__A2 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout319_A net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08986__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09074_ net1226 team_03_WB.instance_to_wrap.core.register_file.registers_state\[173\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[141\] net962 net918
+ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11990__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ net742 _03963_ _03964_ _03965_ _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__o32a_1
XFILLER_0_13_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1130_A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold720 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\] vssd1
+ vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 team_03_WB.instance_to_wrap.core.register_file.registers_state\[566\] vssd1
+ vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold742 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\] vssd1
+ vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10093__C _05811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold753 team_03_WB.instance_to_wrap.core.register_file.registers_state\[131\] vssd1
+ vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 team_03_WB.instance_to_wrap.core.register_file.registers_state\[760\] vssd1
+ vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 team_03_WB.instance_to_wrap.core.register_file.registers_state\[360\] vssd1
+ vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\] vssd1
+ vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold797 team_03_WB.instance_to_wrap.core.register_file.registers_state\[505\] vssd1
+ vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07410__A1 _03351_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _02888_ net2140 net293 vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07961__A2 _03900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ net1049 team_03_WB.instance_to_wrap.core.register_file.registers_state\[203\]
+ net1004 team_03_WB.instance_to_wrap.core.register_file.registers_state\[235\] net922
+ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout855_A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08858_ net861 _04799_ _04796_ net865 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07809_ net1181 team_03_WB.instance_to_wrap.core.register_file.registers_state\[491\]
+ net878 _03750_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08789_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[930\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[898\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[770\]
+ net974 net1070 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10820_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[26\] net307 _06424_ net692
+ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10751_ net527 _06367_ _06368_ net532 net1794 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_98_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08674__B1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10481__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ net1393 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_27_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10682_ net600 _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ net1275 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15140_ net1521 vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ net1408 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ _06613_ net2830 net409 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15071_ net1452 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12283_ net1362 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14022_ clknet_leaf_78_wb_clk_i _01786_ _00387_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[376\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11234_ net1038 _06449_ net650 net701 vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__or4_4
XFILLER_0_120_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ net621 _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ _05947_ _05957_ _05958_ _05959_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__o31ai_1
X_11096_ _06624_ net2823 net424 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output238_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08588__S0 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10047_ net9 net1032 net906 net2547 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__o22a_1
X_14924_ clknet_leaf_126_wb_clk_i _02679_ _01289_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10839__A2 _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__B1 team_03_WB.instance_to_wrap.core.decoder.inst\[31\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 team_03_WB.instance_to_wrap.core.register_file.registers_state\[963\] vssd1
+ vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08362__C1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08901__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\] vssd1
+ vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
X_14855_ clknet_leaf_42_wb_clk_i net1898 _01220_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13806_ clknet_leaf_71_wb_clk_i _01570_ _00171_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[160\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14786_ clknet_leaf_56_wb_clk_i _02550_ _01151_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11998_ _06755_ net469 net450 net2522 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__a22o_1
XANTENNA__07468__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13737_ clknet_leaf_77_wb_clk_i _01501_ _00102_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11264__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ net269 net2483 net522 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13668_ clknet_leaf_13_wb_clk_i _01432_ _00033_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08417__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12619_ net1253 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XANTENNA__11016__A2 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ net1336 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08968__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07928__C1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout507 net509 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_4
X_09830_ net579 _04711_ net543 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o21ai_1
Xfanout518 net520 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_4
Xfanout529 _02923_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
X_09761_ _05654_ _04536_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__and2b_1
X_06973_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[709\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[741\] net729
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a221o_1
XANTENNA__08111__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08712_ _04652_ _04653_ net852 vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__o21a_1
X_09692_ _05276_ _05279_ _05207_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08643_ net1048 team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\] net1003 net940
+ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__o221a_1
XANTENNA__07950__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A _06532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08574_ net1057 _04513_ _04514_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14038__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07459__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07525_ net1095 team_03_WB.instance_to_wrap.core.register_file.registers_state\[582\]
+ net792 team_03_WB.instance_to_wrap.core.register_file.registers_state\[614\] net746
+ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1080_A net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1178_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[245\]
+ net889 vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__or3_1
XFILLER_0_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11007__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout603_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[447\] net768
+ _02869_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1345_A net1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09126_ net849 _05055_ _05067_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__o21ai_4
XANTENNA__09081__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11963__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ net1052 team_03_WB.instance_to_wrap.core.register_file.registers_state\[719\]
+ net1006 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\] net926
+ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ net1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[881\]
+ net894 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or3_1
Xhold550 team_03_WB.instance_to_wrap.CPU_DAT_I\[26\] vssd1 vssd1 vccd1 vccd1 net2134
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout972_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 team_03_WB.instance_to_wrap.core.register_file.registers_state\[232\] vssd1
+ vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\] vssd1
+ vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 team_03_WB.instance_to_wrap.core.register_file.registers_state\[368\] vssd1
+ vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 team_03_WB.instance_to_wrap.core.register_file.registers_state\[276\] vssd1
+ vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__B2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _03600_ net662 vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15146__1527 vssd1 vssd1 vccd1 vccd1 _15146__1527/HI net1527 sky130_fd_sc_hd__conb_1
X_12970_ net1250 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XANTENNA__07147__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08729__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 team_03_WB.instance_to_wrap.core.register_file.registers_state\[76\] vssd1
+ vssd1 vccd1 vccd1 net2834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\] vssd1
+ vssd1 vccd1 vccd1 net2845 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09414__A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _06469_ net2846 net373 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1272 team_03_WB.instance_to_wrap.core.register_file.registers_state\[735\] vssd1
+ vssd1 vccd1 vccd1 net2856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 team_03_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2867
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 net2878
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14640_ clknet_leaf_80_wb_clk_i _02404_ _01005_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\]
+ sky130_fd_sc_hd__dfstp_1
X_11852_ net301 net2026 net381 vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _02798_ _05866_ net320 _06404_ net692 vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__o41a_2
XFILLER_0_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ clknet_leaf_37_wb_clk_i _02335_ _00936_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11246__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ net2124 _06616_ net333 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07869__A net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ net1273 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
X_10734_ team_03_WB.instance_to_wrap.core.pc.current_pc\[14\] _05822_ net601 vssd1
+ vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13453_ net1392 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10665_ team_03_WB.instance_to_wrap.core.ru.state\[3\] team_03_WB.instance_to_wrap.core.ru.state\[4\]
+ team_03_WB.instance_to_wrap.core.ru.state\[5\] vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ net1320 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13384_ net1314 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10596_ team_03_WB.instance_to_wrap.core.ru.state\[4\] _06281_ vssd1 vssd1 vccd1
+ vccd1 _06304_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11954__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15123_ net1504 vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_2
XANTENNA__14800__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12335_ net1407 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054_ net1435 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
X_12266_ net1256 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11706__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ clknet_leaf_88_wb_clk_i _01769_ _00370_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[359\]
+ sky130_fd_sc_hd__dfrtp_1
X_11217_ net271 net2152 net490 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__mux2_1
X_12197_ net1619 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07925__A2 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ _06453_ net703 net695 vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__and3_2
X_11079_ _06617_ net2443 net423 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__mux2_1
XANTENNA__06948__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09324__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ clknet_leaf_39_wb_clk_i _00001_ _01272_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07689__A1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11485__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11065__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A3 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14838_ clknet_leaf_61_wb_clk_i net2273 _01203_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14769_ clknet_leaf_38_wb_clk_i _02533_ _01134_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.READ_I
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08638__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08882__B _04807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07310_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[797\] net800
+ _03246_ net1109 vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08290_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1015\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[983\]
+ net956 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ net1097 team_03_WB.instance_to_wrap.core.register_file.registers_state\[744\]
+ net896 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__or3_1
XANTENNA__07861__A1 net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07172_ net1165 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\]
+ net754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\] net737
+ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__o221a_1
XANTENNA__09063__B1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__C net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__B1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__C1 net1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__A3 net461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout304 _05945_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
Xfanout326 _04833_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
X_09813_ net327 _05545_ _05650_ _05073_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__a22o_1
Xfanout337 net340 vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_8
Xfanout348 net352 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_6
Xfanout359 _04776_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__A1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net358 _05523_ _05678_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a211o_4
X_06956_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[197\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\] net729
+ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a221o_1
XANTENNA__09234__A _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _03391_ _04119_ net539 _02804_ net1088 vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__o32a_1
XANTENNA__11476__A2 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_A net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06887_ _02792_ net1012 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nor2_4
XFILLER_0_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1295_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[6\] net1003
+ net922 _04567_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10099__B net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_A _02863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08629__B1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08557_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[478\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[510\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout818_A net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07508_ _03446_ _03449_ net814 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o21a_1
XANTENNA__07301__A0 _03241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08284__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08488_ net865 _04429_ _04424_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07852__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07439_ net801 _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10450_ team_03_WB.instance_to_wrap.core.pc.current_pc\[4\] team_03_WB.instance_to_wrap.core.pc.current_pc\[3\]
+ team_03_WB.instance_to_wrap.core.pc.current_pc\[2\] team_03_WB.instance_to_wrap.core.pc.current_pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11936__A0 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[462\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[494\] net1069
+ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a221o_1
XANTENNA__08016__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07604__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10381_ _06209_ _06210_ team_03_WB.instance_to_wrap.core.pc.current_pc\[19\] net677
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08801__B1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ net1702 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12051_ _06620_ net2863 net361 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__mux2_1
Xhold380 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\] vssd1
+ vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11377__C net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\] vssd1
+ vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ net2486 net426 _06573_ net519 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XANTENNA__08565__C1 net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14203__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09109__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10911__A1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 _04083_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__buf_4
Xfanout871 _04081_ vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_8
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08317__C1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11393__B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net1357 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
XANTENNA__11467__A2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1080 team_03_WB.instance_to_wrap.core.register_file.registers_state\[324\] vssd1
+ vssd1 vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 team_03_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1 net2675
+ sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net638 _06713_ net478 net379 net2208 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a32o_1
XANTENNA__08963__S0 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12884_ net1322 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14623_ clknet_leaf_109_wb_clk_i _02387_ _00988_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\]
+ sky130_fd_sc_hd__dfstp_1
X_11835_ _06673_ net476 net329 net1923 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07599__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08096__A1 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ clknet_leaf_6_wb_clk_i _02318_ _00919_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[908\]
+ sky130_fd_sc_hd__dfrtp_1
X_11766_ _06597_ net480 net338 net2679 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09832__A2 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ net1390 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10717_ net525 _06348_ _06349_ net530 team_03_WB.instance_to_wrap.ADR_I\[22\] vssd1
+ vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a32o_1
X_14485_ clknet_leaf_72_wb_clk_i _02249_ _00850_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[839\]
+ sky130_fd_sc_hd__dfrtp_1
X_11697_ _06739_ net388 net347 net2084 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08207__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13436_ net1308 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09045__B1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] team_03_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ net841 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09596__A1 _04778_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13367_ net1285 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
X_10579_ net1884 net535 net596 _05889_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a22o_1
XANTENNA__10753__A net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15106_ net1487 vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_2
X_12318_ net1384 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XANTENNA__09319__A _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ net1330 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15037_ clknet_leaf_61_wb_clk_i _02757_ _01402_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__dfrtp_1
X_12249_ net1353 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__inv_2
XANTENNA__11287__C net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07359__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__A2 _05735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08556__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__A1 net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10899__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07790_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[939\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[779\]
+ net770 net1121 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux4_1
XANTENNA__12104__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__S net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09054__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ _05400_ _05401_ net563 vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07531__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ net864 _04352_ _04347_ net848 vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _05321_ _05324_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08342_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\] net917
+ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__o221a_1
XANTENNA__08087__A1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13304__A net1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__B _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08273_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\]
+ net969 team_03_WB.instance_to_wrap.core.register_file.registers_state\[119\] net920
+ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__o221a_1
XANTENNA__07834__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09928__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[818\] net753
+ net1037 _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15145__1526 vssd1 vssd1 vccd1 vccd1 _15145__1526/HI net1526 sky130_fd_sc_hd__conb_1
XFILLER_0_6_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07155_ net1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[416\]
+ net879 _02870_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout301_A _06442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10197__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A _02791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07086_ net1182 net876 team_03_WB.instance_to_wrap.core.register_file.registers_state\[641\]
+ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1210_A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08547__C1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11697__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout670_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10602__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07988_ net1128 _03926_ _03927_ _03929_ net1114 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__a311o_1
XFILLER_0_57_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07770__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ _04150_ _04269_ _04326_ _04386_ net565 net561 vssd1 vssd1 vccd1 vccd1 _05669_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11449__A2 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06939_ _02877_ _02878_ _02880_ _02879_ net744 net808 vssd1 vssd1 vccd1 vccd1 _02881_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11143__C_N net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09511__A1 _05371_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__A0 team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _05089_ _05098_ net562 vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ net870 _04549_ _04550_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a21o_1
XANTENNA__11941__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09589_ _02783_ _02804_ net539 _05528_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__o221a_1
XANTENNA__11433__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _06694_ net386 net353 net2321 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA__13214__A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11551_ net2095 net487 _06790_ net503 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__a22o_1
XANTENNA__11621__A2 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ net129 net1027 net903 net1932 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14270_ clknet_leaf_49_wb_clk_i _02034_ _00635_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[624\]
+ sky130_fd_sc_hd__dfrtp_1
X_11482_ net2558 net399 _06775_ net511 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XANTENNA__11909__A0 _06609_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13221_ net1271 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XANTENNA__07038__C1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10433_ net284 _06251_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__nand3_1
XFILLER_0_85_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07589__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08786__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net1407 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XANTENNA_input64_A gpio_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09139__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ net2877 net676 _06194_ _06196_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__08250__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12103_ net632 _06677_ net469 net445 net2042 vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a32o_1
X_13083_ net1360 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
X_10295_ team_03_WB.instance_to_wrap.core.pc.current_pc\[8\] _06136_ vssd1 vssd1 vccd1
+ vccd1 _06137_ sky130_fd_sc_hd__and2_1
XANTENNA__11137__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14719__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07882__A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__C1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ net632 _06603_ net469 net368 net2285 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__a32o_1
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11688__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10896__B1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07093__S net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 net691 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_4
X_13985_ clknet_leaf_0_wb_clk_i _01749_ _00350_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12101__A3 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12936_ net1293 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XANTENNA__10112__A2 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07513__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12867_ net1296 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13124__A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14606_ clknet_leaf_68_wb_clk_i _02370_ _00971_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_16_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13893__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ _06647_ net466 net329 net2214 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__a22o_1
XANTENNA__08069__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11570__C net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12798_ net1384 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
X_14537_ clknet_leaf_60_wb_clk_i _02301_ _00902_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07277__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07816__A1 net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ net652 _06572_ net464 net337 net2113 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a32o_1
XFILLER_0_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11612__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07816__B2 net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12963__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468_ clknet_leaf_16_wb_clk_i _02232_ _00833_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14249__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ net1423 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XANTENNA__09569__B2 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14399_ clknet_leaf_109_wb_clk_i _02163_ _00764_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11376__A1 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__C1 net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__A1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07675__S0 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08960_ net861 _04898_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11128__B2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[847\]
+ net1149 vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__a21o_1
XANTENNA__11679__A2 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ net581 _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07201__C1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11518__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\] net725
+ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07773_ net1118 _03711_ _03712_ _03714_ net817 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__o311ai_2
XANTENNA__10639__A0 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _05435_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07504__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09443_ _05378_ _05384_ net581 vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout349_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13034__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _05143_ _05159_ _03823_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ net847 _04266_ _04251_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07807__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout516_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1258_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09658__S net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[690\] net913
+ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08480__A1 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06871__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07207_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[434\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[402\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[306\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[274\]
+ net753 net1116 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08187_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[339\]
+ net947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[371\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1425_A net1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07138_ net1158 _03078_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__nand3_1
XANTENNA__11906__A3 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__A2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11001__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07069_ _03008_ _03010_ net805 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__o21a_1
Xoutput260 net260 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
X_10080_ _02925_ _02927_ _05918_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21a_1
XANTENNA__10840__B _05842_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08310__B net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__C1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13770_ clknet_leaf_3_wb_clk_i _01534_ _00135_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net1240 _06449_ net627 net701 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__or4_2
XFILLER_0_35_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12721_ net1311 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net1301 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_307 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _06536_ net2751 net454 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ net1405 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ clknet_leaf_104_wb_clk_i _02086_ _00687_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\]
+ sky130_fd_sc_hd__dfrtp_1
X_11534_ _06434_ net640 net708 net698 vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08471__A1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08472__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ clknet_leaf_105_wb_clk_i _02017_ _00618_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[607\]
+ sky130_fd_sc_hd__dfrtp_1
X_11465_ net2324 net398 _06768_ net502 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11358__A1 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13204_ net1324 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XANTENNA__14541__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10416_ _06008_ _06066_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__and2_1
X_14184_ clknet_leaf_34_wb_clk_i _01948_ _00549_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ net516 net642 _06750_ net408 net2418 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a32o_1
XANTENNA__09420__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ net1391 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
X_10347_ team_03_WB.instance_to_wrap.core.pc.current_pc\[25\] _06182_ net676 vssd1
+ vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07982__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13066_ net1256 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
X_10278_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__inv_2
Xfanout1430 net1431 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__buf_2
X_12017_ _06765_ net463 net365 net2734 vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_14 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__B2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__C1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A3 _06479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12958__A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144__1525 vssd1 vssd1 vccd1 vccd1 _15144__1525/HI net1525 sky130_fd_sc_hd__conb_1
XFILLER_0_75_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13968_ clknet_leaf_81_wb_clk_i _01732_ _00333_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12919_ net1413 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
X_13899_ clknet_leaf_18_wb_clk_i _01663_ _00264_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11833__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08110_ net1086 net892 team_03_WB.instance_to_wrap.core.register_file.registers_state\[538\]
+ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o21a_1
XANTENNA__11801__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08998__C1 net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[557\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[525\]
+ net963 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08462__A1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08041_ _02847_ _03972_ _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold902 team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\] vssd1
+ vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11102__A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\] vssd1
+ vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08214__A1 net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12010__A2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13789__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 team_03_WB.instance_to_wrap.core.register_file.registers_state\[707\] vssd1
+ vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 team_03_WB.instance_to_wrap.core.register_file.registers_state\[691\] vssd1
+ vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\] vssd1
+ vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold957 team_03_WB.instance_to_wrap.core.register_file.registers_state\[677\] vssd1
+ vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07422__C1 net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold968 team_03_WB.instance_to_wrap.core.register_file.registers_state\[771\] vssd1
+ vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _05877_ net1878 net287 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold979 team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\] vssd1
+ vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10572__A2 net537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08943_ net1045 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\]
+ net999 team_03_WB.instance_to_wrap.core.register_file.registers_state\[619\] net939
+ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout299_A _06495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A1 _05073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08874_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07725__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1006_A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07027__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07825_ net807 _03765_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__and3_1
XANTENNA__11194__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout466_A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07756_ net1118 _03693_ _03694_ _03696_ net1108 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__a311o_1
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06866__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10088__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__A _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07489__C1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ _03624_ _03628_ net1138 vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08150__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1375_A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ net578 _05354_ _05367_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09357_ _04984_ _05297_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11711__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08308_ net1217 _04248_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__o21a_1
XANTENNA__07697__A team_03_WB.instance_to_wrap.core.decoder.inst\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08292__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11052__A3 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _04646_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[50\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\]
+ net948 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11250_ net516 net635 _06692_ net415 net2348 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a32o_1
XANTENNA__08205__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09402__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10201_ _02990_ _06041_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07413__C1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11181_ net694 net712 net296 vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10563__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _04354_ _02770_ net671 vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08321__A net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14940_ clknet_leaf_40_wb_clk_i _02695_ _01305_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09136__B _05076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ net2 net1033 net907 net2873 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o22a_1
XANTENNA__11385__C net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07716__B1 net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ clknet_leaf_38_wb_clk_i _02635_ _01236_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.prev_busy
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A3 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13822_ clknet_leaf_48_wb_clk_i _01586_ _00187_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[176\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14094__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09564__S0 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13753_ clknet_leaf_93_wb_clk_i _01517_ _00118_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10965_ net830 _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12704_ net1408 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ clknet_leaf_91_wb_clk_i _01448_ _00049_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08692__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10896_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[14\] net308 net685 vssd1
+ vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a21o_1
XANTENNA__08692__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11028__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ net1364 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ net1338 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09641__B1 _05582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07400__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11517_ _06631_ net2492 net395 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
X_14305_ clknet_leaf_129_wb_clk_i _02069_ _00670_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07652__C1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ net1304 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold209 net194 vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
X_14236_ clknet_leaf_126_wb_clk_i _02000_ _00601_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\]
+ sky130_fd_sc_hd__dfrtp_1
X_11448_ _06434_ net640 net708 net825 vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11200__A0 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14167_ clknet_leaf_87_wb_clk_i _01931_ _00532_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[521\]
+ sky130_fd_sc_hd__dfrtp_1
X_11379_ net712 _06518_ net697 vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ net1413 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
X_14098_ clknet_leaf_102_wb_clk_i _01862_ _00463_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08231__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ net1355 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
XANTENNA__11295__C net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__buf_2
Xfanout1271 net1277 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_4
XFILLER_0_20_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14437__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1282 net1283 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__buf_2
Xfanout1293 net1294 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_2
X_07610_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[985\]
+ net783 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1017\] net1159
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__o221a_1
X_08590_ net846 _04518_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o21ba_4
XANTENNA__08377__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07541_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[486\]
+ net877 _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14587__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07472_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[693\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\] net762 net726
+ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09211_ net605 _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10936__A team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09142_ _04149_ _04208_ net552 vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__B1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[45\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[13\]
+ net964 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09181__A1_N net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__S net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08024_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[177\]
+ net887 net1117 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold710 team_03_WB.instance_to_wrap.core.register_file.registers_state\[762\] vssd1
+ vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\] vssd1
+ vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_03_WB.instance_to_wrap.ADR_I\[5\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold743 team_03_WB.instance_to_wrap.core.register_file.registers_state\[125\] vssd1
+ vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[602\] vssd1
+ vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 team_03_WB.instance_to_wrap.core.register_file.registers_state\[463\] vssd1
+ vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__A1 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 team_03_WB.instance_to_wrap.core.register_file.registers_state\[556\] vssd1
+ vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\] vssd1
+ vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11486__B net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09975_ _02921_ net1822 net295 vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__mux2_1
XANTENNA__07683__C net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\] vssd1
+ vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08141__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08926_ net1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[75\]
+ net998 team_03_WB.instance_to_wrap.core.register_file.registers_state\[107\] net940
+ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09699__B1 net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07980__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _04797_ _04798_ net941 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__mux2_1
XANTENNA__09794__S0 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07808_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[459\]
+ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__and2_1
XANTENNA__10610__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08788_ _04728_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__and2_1
XANTENNA__07191__S net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11258__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ _03669_ _03677_ net614 _03660_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o211a_2
XFILLER_0_71_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10549__C _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ _05730_ net602 vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08674__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09871__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09409_ net552 _04985_ _04180_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13954__CLK clknet_leaf_129_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10481__B2 net2345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ net317 _06314_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ net1303 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11430__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12351_ net1377 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_67_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11302_ _06612_ net2596 net409 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__mux2_1
X_15143__1524 vssd1 vssd1 vccd1 vccd1 _15143__1524/HI net1524 sky130_fd_sc_hd__conb_1
X_15070_ net1451 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12282_ net1371 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ clknet_leaf_108_wb_clk_i _01785_ _00386_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[375\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ net266 net2260 net493 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10536__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__A1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__S net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ net694 net709 net299 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__or3b_1
XANTENNA__08051__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ net679 net284 team_03_WB.instance_to_wrap.core.pc.current_pc\[1\] vssd1 vssd1
+ vccd1 vccd1 _05959_ sky130_fd_sc_hd__a21bo_1
X_11095_ net828 net271 vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08588__S1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ net10 net1035 net908 net2675 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
X_14923_ clknet_leaf_126_wb_clk_i _02678_ _01288_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07165__A1 _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[12\] vssd1 vssd1 vccd1
+ vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1006\] vssd1
+ vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_03_WB.instance_to_wrap.CPU_DAT_I\[5\] vssd1 vssd1 vccd1 vccd1 net1676
+ sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ clknet_leaf_41_wb_clk_i net1968 _01219_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ clknet_leaf_105_wb_clk_i _01569_ _00170_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[159\]
+ sky130_fd_sc_hd__dfrtp_1
X_14785_ clknet_leaf_41_wb_clk_i _02549_ _01150_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11997_ net297 net2474 net451 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13736_ clknet_leaf_26_wb_clk_i _01500_ _00101_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ _06529_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11264__A3 _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09610__A _05551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13667_ clknet_leaf_19_wb_clk_i _01431_ _00032_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10879_ net313 net311 net322 _02779_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08417__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ net1249 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09614__B1 net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ net1278 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12549_ net1275 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06979__A1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14219_ clknet_leaf_36_wb_clk_i _01983_ _00584_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[573\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15199_ net1574 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_65_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10527__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A1 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__B1 net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09760_ _04777_ _05072_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__a21bo_1
X_06972_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[581\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[613\] net743
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a221o_1
X_08711_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[132\]
+ net975 team_03_WB.instance_to_wrap.core.register_file.registers_state\[164\] net939
+ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__o221a_1
X_09691_ _05623_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1090 net1092 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__buf_2
X_08642_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\]
+ net979 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08573_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[445\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[413\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[317\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\]
+ net967 net1069 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08105__B1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07524_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[678\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[646\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07455_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[85\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[117\] net726
+ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06863__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1073_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07386_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[415\] net791
+ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__or2_1
XANTENNA__11412__A0 _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09125_ net1077 _05060_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09081__A1 net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1240_A net1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11963__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1338_A net1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07975__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _04992_ _04997_ net871 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ net1089 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1009\]
+ net893 _03948_ net1146 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__o311a_1
XANTENNA__14602__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\] vssd1
+ vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10605__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold551 team_03_WB.instance_to_wrap.ADR_I\[3\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10518__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__A1 _06422_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 team_03_WB.instance_to_wrap.core.register_file.registers_state\[279\] vssd1
+ vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold573 team_03_WB.instance_to_wrap.core.register_file.registers_state\[811\] vssd1
+ vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 team_03_WB.instance_to_wrap.core.register_file.registers_state\[411\] vssd1
+ vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold595 team_03_WB.instance_to_wrap.core.register_file.registers_state\[248\] vssd1
+ vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11191__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _05883_ net1861 net293 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08909_ net1043 team_03_WB.instance_to_wrap.core.register_file.registers_state\[652\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[684\] net917
+ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a221o_1
XANTENNA__11479__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ net326 _05449_ _05513_ _05436_ _05830_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1240 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\] vssd1
+ vssd1 vccd1 vccd1 net2824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1251 team_03_WB.instance_to_wrap.core.register_file.registers_state\[222\] vssd1
+ vssd1 vccd1 vccd1 net2835 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10151__A0 _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ _06454_ net2809 net373 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__mux2_1
Xhold1262 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\] vssd1
+ vssd1 vccd1 vccd1 net2846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 team_03_WB.instance_to_wrap.core.register_file.registers_state\[723\] vssd1
+ vssd1 vccd1 vccd1 net2857 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1284 team_03_WB.instance_to_wrap.wb.curr_state\[1\] vssd1 vssd1 vccd1 vccd1 net2868
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08895__B2 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1295 team_03_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1 net2879
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11851_ net302 net2146 net382 vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__mux2_1
XANTENNA__09133__C net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10802_ net314 net312 net323 _02778_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14570_ clknet_leaf_2_wb_clk_i _02334_ _00935_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[924\]
+ sky130_fd_sc_hd__dfrtp_1
X_11782_ net2633 _06615_ net332 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10733_ net2428 net530 net528 _06358_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13521_ net1281 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07855__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ net1393 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ team_03_WB.instance_to_wrap.core.ru.state\[4\] team_03_WB.instance_to_wrap.core.ru.state\[5\]
+ team_03_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__o21a_1
XANTENNA_input94_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07588__C net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10206__A1 _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11403__A0 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_775 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12403_ net1267 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XANTENNA__07607__C1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13383_ net1423 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XANTENNA__09072__A1 _03105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10595_ net1134 net1899 net842 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11954__A1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15122_ net1503 vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_2
X_12334_ net1338 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XANTENNA__14282__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15053_ net1434 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
X_12265_ net1252 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10509__A2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ clknet_leaf_92_wb_clk_i _01768_ _00369_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[358\]
+ sky130_fd_sc_hd__dfrtp_1
X_11216_ net300 net2690 net493 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08032__C1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12196_ net1586 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ net502 net651 _06650_ net418 net1960 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a32o_1
XFILLER_0_78_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11078_ net829 net275 vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and2_2
XANTENNA__06948__B _02889_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ team_03_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _05905_ sky130_fd_sc_hd__nand2_1
X_14906_ clknet_leaf_37_wb_clk_i _00000_ _01271_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.ru.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07125__A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__B2 _06332_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14837_ clknet_leaf_32_wb_clk_i net2038 _01202_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11890__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09043__C _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08638__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14768_ clknet_leaf_37_wb_clk_i _02532_ _01133_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.i_hit
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13719_ clknet_leaf_73_wb_clk_i _01483_ _00084_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11642__B1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14699_ clknet_leaf_53_wb_clk_i _02463_ _01064_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11081__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07240_ net1185 team_03_WB.instance_to_wrap.core.register_file.registers_state\[968\]
+ net774 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\] net1148
+ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07171_ net1163 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\]
+ net754 team_03_WB.instance_to_wrap.core.register_file.registers_state\[115\] net724
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__o221a_1
XANTENNA__09063__A1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11945__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07074__B1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08271__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14775__CLK clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11110__A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _05925_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07377__A1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07916__A3 net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ net575 _04957_ _05753_ _04777_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__o211a_1
Xfanout327 _04833_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_8
Xfanout349 net351 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_6
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06955_ net1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[69\]
+ net790 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\] net744
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a221o_1
X_09743_ _05073_ _05601_ _05682_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a211o_1
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout281_A _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ _05614_ _05615_ net359 vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__o21a_1
X_06886_ _02823_ _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__or2_1
XANTENNA__08877__B2 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08625_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\] net979
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or2_1
X_15142__1523 vssd1 vssd1 vccd1 vccd1 _15142__1523/HI net1523 sky130_fd_sc_hd__conb_1
XANTENNA__11881__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08629__A1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08556_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[350\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[382\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06874__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10436__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ net810 _03447_ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11633__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _04425_ _04426_ _04428_ _04427_ net926 net862 vssd1 vssd1 vccd1 vccd1 _04429_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout713_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07438_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[212\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[244\] net742
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ net1106 _03309_ _03310_ _03304_ _03305_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13500__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[334\]
+ net995 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\] net1203
+ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10380_ net283 _06145_ _06206_ net677 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__o31a_1
XANTENNA__08801__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__B net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09039_ _04977_ _04978_ _04979_ _04980_ net862 net944 vssd1 vssd1 vccd1 vccd1 _04981_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11020__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12050_ _06619_ net2785 net361 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__mux2_1
Xhold370 _02588_ vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold381 net103 vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07368__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ net276 net657 net707 net825 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__and4_1
Xhold392 team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\] vssd1
+ vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10911__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout850 net851 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_4
Xfanout861 net862 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout883 net884 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_2
XANTENNA__08317__B1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout894 net901 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08868__A1 _02937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11393__C net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ net1368 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 team_03_WB.instance_to_wrap.core.register_file.registers_state\[323\] vssd1
+ vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 team_03_WB.instance_to_wrap.core.register_file.registers_state\[815\] vssd1
+ vssd1 vccd1 vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1092 team_03_WB.instance_to_wrap.core.register_file.registers_state\[635\] vssd1
+ vssd1 vccd1 vccd1 net2676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11903_ net636 _06712_ net475 net379 net2255 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__a32o_1
XANTENNA__11872__A0 _06545_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08963__S1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12786__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12883_ net1259 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14622_ clknet_leaf_57_wb_clk_i _02386_ _00987_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_16_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11834_ _06672_ net478 net330 net2164 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10427__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14648__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__B1 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14553_ clknet_leaf_111_wb_clk_i _02317_ _00918_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[907\]
+ sky130_fd_sc_hd__dfrtp_1
X_11765_ net650 _06595_ net459 net337 net2027 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_82_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09832__A3 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10716_ _05842_ net601 vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nand2_1
X_13504_ net1391 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11696_ _06738_ net386 net345 net1941 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__a22o_1
X_14484_ clknet_leaf_91_wb_clk_i _02248_ _00849_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[838\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08207__C _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13435_ net1400 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10647_ team_03_WB.instance_to_wrap.core.decoder.inst\[14\] team_03_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ net840 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07111__C net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08253__C1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ net1291 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
X_10578_ net1774 net534 net595 _05888_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08504__A _04080_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ net1486 vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_2
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12317_ net1382 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
X_13297_ net1392 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15036_ clknet_leaf_61_wb_clk_i _02756_ _01401_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__dfrtp_1
X_12248_ net1362 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08556__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12179_ net1661 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14178__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11863__B1 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08410_ _04348_ _04349_ _04351_ _04350_ net943 net861 vssd1 vssd1 vccd1 vccd1 _04352_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11804__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09390_ _05323_ _05327_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__or2_1
XANTENNA__09808__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10418__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ net935 _04281_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11615__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10969__A2 _05082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08272_ _04212_ _04213_ net859 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07302__B _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08492__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07223_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[786\] net787
+ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ _03093_ _03095_ net1112 vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10663__B net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11394__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06860__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07085_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[513\] net792
+ net731 _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09944__S net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ net1100 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\]
+ net900 _03928_ net1147 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__o311a_1
XFILLER_0_138_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout663_A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07770__A1 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06938_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[612\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[580\]
+ net769 vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__mux2_1
X_09726_ net358 _05438_ _05665_ _04820_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__a221o_1
XANTENNA__11854__A0 _06453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _05293_ _05298_ _05597_ _05294_ _05285_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a311oi_4
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout830_A _06387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _02811_ sky130_fd_sc_hd__nand3b_4
XANTENNA_fanout928_A _04088_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11714__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08608_ net864 _04541_ _04544_ net843 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__a31o_1
X_09588_ _04071_ _04382_ net663 _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a22o_1
XANTENNA__11941__C _06562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11606__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08539_ net1056 _04479_ _04480_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11015__A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net651 _06660_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07286__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10501_ net2472 net1028 net903 net2316 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08027__C net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09027__A1 net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ net637 net706 _06541_ net824 vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__and4_1
XFILLER_0_68_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ net1309 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10432_ _06020_ _06022_ _06061_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or3_1
XANTENNA__07038__B1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12031__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08786__B1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ net1376 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ net283 _06147_ _06195_ net676 vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__o31a_1
X_12102_ _06797_ net478 net445 net2010 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ net1365 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10294_ team_03_WB.instance_to_wrap.core.pc.current_pc\[7\] team_03_WB.instance_to_wrap.core.pc.current_pc\[6\]
+ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__and3_1
XANTENNA_input57_A gpio_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__A2 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12033_ _06774_ net479 net367 net2673 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14320__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_2
XFILLER_0_75_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12098__B1 net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_4
X_13984_ clknet_leaf_134_wb_clk_i _01748_ _00349_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__A0 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__A1 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12935_ net1399 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07513__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08710__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12866_ net1364 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ clknet_leaf_106_wb_clk_i _02369_ _00970_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[959\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11817_ _06645_ net473 net330 net1944 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a22o_1
XANTENNA__11570__D net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797_ net1372 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07277__B1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ clknet_leaf_34_wb_clk_i _02300_ _00901_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[890\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _06571_ net481 net339 net2289 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09018__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__A1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[26\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09018__B2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14467_ clknet_leaf_26_wb_clk_i _02231_ _00832_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ _06721_ net387 net344 net1942 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13140__A net1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13418_ net1308 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XANTENNA__09569__A2 _04235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12022__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__C1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14398_ clknet_leaf_48_wb_clk_i _02162_ _00763_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[752\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08234__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08777__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ net1294 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15141__1522 vssd1 vssd1 vccd1 vccd1 _15141__1522/HI net1522 sky130_fd_sc_hd__conb_1
XANTENNA__07675__S1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11128__A2 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15019_ clknet_leaf_62_wb_clk_i _02739_ _01384_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__dfrtp_1
X_07910_ net1159 _03845_ _03846_ _03848_ _03851_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08890_ net585 _04830_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07841_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[586\]
+ net787 team_03_WB.instance_to_wrap.core.register_file.registers_state\[618\] net738
+ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12089__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ net1108 _03704_ _03705_ _03713_ net1143 vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__a311o_1
XFILLER_0_100_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06960__C1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ _05371_ _05438_ _05450_ _05452_ _05448_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__a221o_2
XFILLER_0_91_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11836__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09442_ _05381_ _05383_ net567 vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__mux2_1
XANTENNA__09512__B _05453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07313__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ _05313_ _05314_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08324_ _04257_ _04260_ _04265_ net864 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08255_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[562\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[530\]
+ net948 vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1153_A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07206_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[466\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[498\] net1142
+ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12013__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08217__C1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ net855 _04124_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08768__B1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07137_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[832\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[864\] net1150
+ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1320_A net1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1418_A net1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__C net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__B1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\] net790
+ net729 _03009_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout780_A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput250 net250 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XANTENNA__07991__A1 _02872_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput261 net261 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XANTENNA_fanout878_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__B2 _02870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07194__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire1014 _02817_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_96_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07743__A1 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08940__B1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _03682_ _05041_ net541 vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11827__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ net1245 net831 vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__nand2_4
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12095__A3 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ net1428 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ net1257 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ net269 net2618 net454 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ net1427 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08456__C1 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10802__A1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ clknet_leaf_94_wb_clk_i _02085_ _00686_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\]
+ sky130_fd_sc_hd__dfrtp_1
X_11533_ net2121 net489 _06784_ net519 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ net651 _06589_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nor2_1
XANTENNA__12004__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ clknet_leaf_6_wb_clk_i _02016_ _00617_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[606\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11358__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ team_03_WB.instance_to_wrap.core.pc.current_pc\[11\] _06139_ team_03_WB.instance_to_wrap.core.pc.current_pc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ net1264 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
X_14183_ clknet_leaf_64_wb_clk_i _01947_ _00548_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[537\]
+ sky130_fd_sc_hd__dfrtp_1
X_11395_ net714 net266 net698 vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07026__A3 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__C net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ _06179_ _06181_ net282 vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__mux2_1
X_13134_ net1340 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XANTENNA__14836__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13710__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13065_ net1255 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
X_10277_ _06115_ _06118_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1420 net1426 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__buf_4
X_12016_ _06764_ net468 net368 net2714 vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a22o_1
Xfanout1431 net1432 vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11530__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14986__CLK clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11818__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ clknet_leaf_97_wb_clk_i _01731_ _00332_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12086__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__A net1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12918_ net1343 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08695__C1 net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ clknet_leaf_3_wb_clk_i _01662_ _00263_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[252\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12849_ net1312 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ clknet_leaf_76_wb_clk_i _02283_ _00884_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[873\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08040_ net816 _03977_ _03979_ _03981_ net720 vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__a41o_1
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold903 team_03_WB.instance_to_wrap.core.register_file.registers_state\[747\] vssd1
+ vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11102__B net270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold914 team_03_WB.instance_to_wrap.core.register_file.registers_state\[625\] vssd1
+ vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10557__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold925 team_03_WB.instance_to_wrap.core.register_file.registers_state\[369\] vssd1
+ vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold936 team_03_WB.instance_to_wrap.core.register_file.registers_state\[229\] vssd1
+ vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[759\] vssd1
+ vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[576\] vssd1
+ vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09991_ _05876_ net2306 net291 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__mux2_1
Xhold969 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\] vssd1
+ vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10941__B _05746_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ _04880_ _04883_ team_03_WB.instance_to_wrap.core.decoder.inst\[18\] vssd1
+ vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08873_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__nor2_1
XANTENNA__07725__A1 net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ net1079 team_03_WB.instance_to_wrap.core.register_file.registers_state\[202\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[234\] net728
+ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09190__A3 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07755_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[428\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[396\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[300\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[268\]
+ net761 net1118 vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12077__A3 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout459_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07489__B1 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _03626_ _03627_ net1152 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__a21o_1
XANTENNA__08139__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08150__A1 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09425_ net565 _05366_ _05359_ net581 vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1270_A net1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout626_A net645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1368_A net1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07978__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14709__CLK clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ _04984_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2_2
XANTENNA__11037__B2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06882__A team_03_WB.instance_to_wrap.core.decoder.inst\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08989__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08307_ net1062 _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07697__B net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ _03208_ _05223_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10608__S net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10796__A0 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__S net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08238_ net552 _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13733__CLK clknet_leaf_108_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[948\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[916\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ _02990_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__nor2_1
XANTENNA__07413__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11180_ net2420 net419 _06670_ net512 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10851__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11760__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _03313_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10062_ net13 net1036 net909 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1
+ vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
X_14870_ clknet_leaf_53_wb_clk_i net2055 _01235_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10720__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ clknet_leaf_67_wb_clk_i _01585_ _00186_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[175\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11276__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13752_ clknet_leaf_12_wb_clk_i _01516_ _00117_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ _06542_ _06543_ _06544_ _06399_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__o211a_4
XFILLER_0_134_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11815__A3 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15140__1521 vssd1 vssd1 vccd1 vccd1 _15140__1521/HI net1521 sky130_fd_sc_hd__conb_1
XANTENNA__08049__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12703_ net1377 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13683_ clknet_leaf_113_wb_clk_i _01447_ _00048_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10895_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[14\] net306 vssd1
+ vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11028__A1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ net1370 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XANTENNA__08483__S net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08444__A2 _04384_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ net1268 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07101__C1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ clknet_leaf_132_wb_clk_i _02068_ _00669_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[658\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07652__B1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ net264 net2762 net396 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12496_ net1418 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
XFILLER_0_48_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ clknet_leaf_29_wb_clk_i _01999_ _00600_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[589\]
+ sky130_fd_sc_hd__dfrtp_1
X_11447_ net2512 net399 _06762_ net519 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10539__B1 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08601__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ clknet_leaf_84_wb_clk_i _01930_ _00531_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[520\]
+ sky130_fd_sc_hd__dfrtp_1
X_11378_ net516 net640 _06741_ net408 net2215 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07955__A1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _06167_ _06166_ net282 vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__mux2_1
X_13117_ net1383 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ clknet_leaf_94_wb_clk_i _01861_ _00462_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ net1363 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12969__A net1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_2
Xfanout1261 net1270 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
Xfanout1272 net1277 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_2
Xfanout1283 net1295 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_4
XANTENNA__06967__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08380__A1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1294 net1295 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_2
XFILLER_0_89_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14999_ clknet_leaf_126_wb_clk_i net47 _01364_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07540_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[454\]
+ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07471_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[533\] net762
+ net741 _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ net438 _05146_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07798__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__B net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ net546 _04208_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nor2_1
XANTENNA__13756__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11113__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ _03105_ _04985_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_86_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08840__C1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08023_ net1081 net887 team_03_WB.instance_to_wrap.core.register_file.registers_state\[145\]
+ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold700 team_03_WB.instance_to_wrap.core.register_file.registers_state\[470\] vssd1
+ vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold711 team_03_WB.instance_to_wrap.core.register_file.registers_state\[926\] vssd1
+ vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 net223 vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold733 team_03_WB.instance_to_wrap.core.register_file.registers_state\[867\] vssd1
+ vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08738__A3 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold744 team_03_WB.instance_to_wrap.core.register_file.registers_state\[675\] vssd1
+ vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07964__C net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 team_03_WB.instance_to_wrap.core.register_file.registers_state\[896\] vssd1
+ vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10671__B _05583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold766 team_03_WB.instance_to_wrap.core.register_file.registers_state\[855\] vssd1
+ vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold777 team_03_WB.instance_to_wrap.core.register_file.registers_state\[746\] vssd1
+ vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10163__S net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold788 team_03_WB.instance_to_wrap.core.register_file.registers_state\[394\] vssd1
+ vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _03488_ net2226 net294 vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__mux2_1
XANTENNA__11486__C net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[426\] vssd1
+ vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08141__B net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1116_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__S net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _04865_ _04866_ net852 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12879__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09699__A1 _04816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[672\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[640\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__mux2_1
XANTENNA__09794__S1 net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11029__C_N net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06877__A _02808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07807_ net1090 team_03_WB.instance_to_wrap.core.register_file.registers_state\[331\]
+ net791 team_03_WB.instance_to_wrap.core.register_file.registers_state\[363\] net1147
+ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_135_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout743_A net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[962\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[994\] net1070
+ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11258__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07738_ net608 _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout910_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07669_ net1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[254\]
+ net885 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13503__A net1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ _05348_ _05349_ net555 vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__mux2_1
X_10680_ _06307_ net530 vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nor2_1
XANTENNA__10481__A2 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _05204_ _05207_ _05279_ _05280_ _05201_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__o311a_2
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11430__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07634__B1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ net1384 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11301_ _06611_ net2841 net409 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__mux2_1
X_12281_ net1353 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__S0 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14020_ clknet_leaf_18_wb_clk_i _01784_ _00385_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[374\]
+ sky130_fd_sc_hd__dfrtp_1
X_11232_ _06550_ net2220 net492 vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07398__C1 net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ net498 net647 _06659_ net417 net1760 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10114_ _05952_ _05953_ _05956_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _06623_ net2775 net422 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__mux2_1
X_10045_ net11 net1036 net908 net2827 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a22o_1
X_14922_ clknet_leaf_125_wb_clk_i _02677_ _01287_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09154__A3 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08898__C1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__A1 net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 team_03_WB.instance_to_wrap.core.register_file.registers_state\[951\] vssd1
+ vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10839__A4 _06403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1000\] vssd1
+ vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\] vssd1
+ vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ clknet_leaf_53_wb_clk_i net2059 _01218_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
Xhold93 _02576_ vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ clknet_leaf_9_wb_clk_i _01568_ _00169_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[158\]
+ sky130_fd_sc_hd__dfrtp_1
X_14784_ clknet_leaf_32_wb_clk_i _02548_ _01149_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10102__A _05925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08114__A1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ _06509_ net2451 net449 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13779__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13735_ clknet_leaf_65_wb_clk_i _01499_ _00100_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10947_ net690 _05757_ _06399_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07873__B1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13666_ clknet_leaf_127_wb_clk_i _01430_ _00031_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10878_ net691 _05632_ net586 vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07411__A net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12617_ net1248 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ net1337 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12548_ net1311 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
XANTENNA__08822__C1 net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__B2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net1356 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14218_ clknet_leaf_10_wb_clk_i _01982_ _00583_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[572\]
+ sky130_fd_sc_hd__dfrtp_1
X_15198_ net911 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__A1 net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11079__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ clknet_leaf_108_wb_clk_i _01913_ _00514_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08050__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout509 net514 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06971_ net1140 _02912_ net718 vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11807__S net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[4\] net1002
+ net923 _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__o211a_1
XANTENNA__09145__A3 _04323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09690_ net582 _05624_ _05625_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a31o_2
XANTENNA__14554__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07156__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1080 net1088 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_4
X_08641_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\]
+ net979 net1073 vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__mux4_1
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06903__A2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08572_ net1228 team_03_WB.instance_to_wrap.core.register_file.registers_state\[477\]
+ net960 team_03_WB.instance_to_wrap.core.register_file.registers_state\[509\] net1202
+ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07523_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[550\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\]
+ net775 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07454_ net739 _03392_ _03393_ _03394_ _03395_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__o32a_1
XFILLER_0_76_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07385_ _03325_ _03326_ net1157 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08136__B _03391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1066_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ net866 _05065_ net844 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09055_ net1062 _04995_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a21o_1
XANTENNA__07092__A1 net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1233_A net1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08006_ net1179 team_03_WB.instance_to_wrap.core.register_file.registers_state\[977\]
+ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09248__A _04294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold530 team_03_WB.instance_to_wrap.core.register_file.registers_state\[366\] vssd1
+ vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08152__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold541 team_03_WB.instance_to_wrap.core.register_file.registers_state\[703\] vssd1
+ vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 net193 vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold563 team_03_WB.instance_to_wrap.core.register_file.registers_state\[915\] vssd1
+ vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold574 team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\] vssd1
+ vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1400_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold585 team_03_WB.instance_to_wrap.core.register_file.registers_state\[487\] vssd1
+ vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 net155 vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ _03844_ _03863_ net661 vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nor3_2
XANTENNA_fanout860_A _04083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11717__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _04848_ _04849_ net1210 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__o21a_1
XANTENNA__11479__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10621__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ net1016 _03109_ _04820_ _05827_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\] vssd1
+ vssd1 vccd1 vccd1 net2814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 team_03_WB.instance_to_wrap.core.register_file.registers_state\[595\] vssd1
+ vssd1 vccd1 vccd1 net2825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1252 team_03_WB.instance_to_wrap.core.register_file.registers_state\[830\] vssd1
+ vssd1 vccd1 vccd1 net2836 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[0\] net1005
+ net925 _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__o211a_1
XANTENNA__13921__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1263 team_03_WB.instance_to_wrap.core.register_file.registers_state\[204\] vssd1
+ vssd1 vccd1 vccd1 net2847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 team_03_WB.instance_to_wrap.core.register_file.registers_state\[140\] vssd1
+ vssd1 vccd1 vccd1 net2858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 team_03_WB.instance_to_wrap.core.register_file.registers_state\[82\] vssd1
+ vssd1 vccd1 vccd1 net2869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11850_ net275 net2143 net383 vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ net280 net2295 net521 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
X_11781_ net2768 _06614_ net334 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13233__A net1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ net1279 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
X_10732_ team_03_WB.instance_to_wrap.core.pc.current_pc\[15\] _05646_ net601 vssd1
+ vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13451_ net1396 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
X_10663_ _06300_ net604 net1137 vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__and3b_1
XANTENNA__09057__C1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12402_ net1389 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
XANTENNA__07607__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13382_ net1308 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
X_10594_ team_03_WB.instance_to_wrap.core.ru.prev_busy team_03_WB.instance_to_wrap.core.ru.state\[3\]
+ _06281_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__and3_1
XANTENNA_input87_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08804__C1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10975__A_N _02829_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14427__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15121_ net1502 vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_2
XFILLER_0_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12333_ net1268 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09158__A net570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ net1584 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12264_ net1284 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ clknet_leaf_111_wb_clk_i _01767_ _00368_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11706__A2 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11215_ _06483_ net2378 net493 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__mux2_1
X_12195_ net1622 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__14577__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ net274 net704 net696 vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__and3_1
XANTENNA__10390__A1 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11077_ _06616_ net2561 net422 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10028_ team_03_WB.instance_to_wrap.wb.curr_state\[1\] net1 vssd1 vssd1 vccd1 vccd1
+ _05904_ sky130_fd_sc_hd__and2_1
X_14905_ clknet_leaf_30_wb_clk_i _00010_ _01270_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09532__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14836_ clknet_leaf_32_wb_clk_i net1988 _01201_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11890__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07840__S net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08099__B1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ clknet_leaf_37_wb_clk_i _02531_ _01132_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.d_hit
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11979_ net303 net2485 net450 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10445__A2 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ clknet_leaf_86_wb_clk_i _01482_ _00083_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14698_ clknet_leaf_53_wb_clk_i _02462_ _01063_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08237__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07310__A2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09048__C1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ clknet_leaf_95_wb_clk_i _01413_ _00014_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07170_ _03110_ _03111_ net737 vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06980__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07074__A1 net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10706__S net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11158__B1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11110__B net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10905__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ net574 _04650_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__nand2_1
Xfanout317 _05387_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
Xfanout328 net331 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_8
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_6
XANTENNA__13944__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09742_ _05527_ _05654_ _05683_ _04777_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__a2bb2o_1
X_06954_ _02894_ _02895_ net729 vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__mux2_1
XANTENNA__08326__A1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06858__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09673_ net576 _05570_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nor2_1
XANTENNA__08877__A2 _04770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06885_ _02808_ _02817_ _02820_ _02826_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_119_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout274_A _06446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08624_ net442 net434 _04565_ net553 vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__o31a_1
XFILLER_0_94_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08555_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[446\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[414\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[318\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[286\]
+ net954 net1066 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout1183_A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout539_A net540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07506_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[199\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\] net733
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1019\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[987\]
+ net988 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ net1162 team_03_WB.instance_to_wrap.core.register_file.registers_state\[84\]
+ net756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[116\] net724
+ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__o221a_1
XANTENNA__10841__C1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1350_A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ net724 _03299_ _03300_ net1138 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ net856 _05047_ _05048_ _05046_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__a31o_1
XFILLER_0_126_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07299_ _03217_ _03224_ _03233_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__10616__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[1008\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\]
+ net982 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11149__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\] vssd1
+ vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 team_03_WB.instance_to_wrap.core.register_file.registers_state\[436\] vssd1
+ vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 net217 vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A1 net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ net502 net651 _06572_ net425 net2177 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a32o_1
Xhold393 team_03_WB.instance_to_wrap.core.register_file.registers_state\[237\] vssd1
+ vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08565__B2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07773__C1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net841 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout851 _04084_ vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
Xfanout862 _04083_ vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_4
Xfanout873 net884 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_4
XANTENNA__08317__A1 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout884 _02845_ vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_4
Xfanout895 net901 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
X_12951_ net1417 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1060 team_03_WB.instance_to_wrap.core.register_file.registers_state\[496\] vssd1
+ vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07525__C1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1071 team_03_WB.instance_to_wrap.core.register_file.registers_state\[91\] vssd1
+ vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_9_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11902_ net630 _06711_ net468 net380 net2520 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__a32o_1
XFILLER_0_119_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1082 team_03_WB.instance_to_wrap.core.register_file.registers_state\[192\] vssd1
+ vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net1420 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
Xhold1093 team_03_WB.instance_to_wrap.core.register_file.registers_state\[730\] vssd1
+ vssd1 vccd1 vccd1 net2677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14621_ clknet_leaf_63_wb_clk_i _02385_ _00986_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[975\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_115_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11833_ _06670_ net476 net329 net2051 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09817__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14552_ clknet_leaf_10_wb_clk_i _02316_ _00917_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07828__B1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11764_ _06594_ net471 net338 net2426 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13503_ net1328 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10715_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] net600 vssd1 vssd1 vccd1
+ vccd1 _06348_ sky130_fd_sc_hd__or2_1
X_14483_ clknet_leaf_113_wb_clk_i _02247_ _00848_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[837\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11695_ _06737_ net386 net345 net2441 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11910__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13817__CLK clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ net1308 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ net1229 net1823 net842 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09045__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11388__B1 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ net1321 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ net1862 net535 net596 _05887_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12307__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08504__B _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ net1485 vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_2
XANTENNA__10060__B1 net909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net1355 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
X_13296_ net1330 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15035_ clknet_leaf_40_wb_clk_i _02755_ _01400_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12247_ net1696 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09753__B1 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09616__A net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ net1616 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13138__A net1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ net1038 net831 net279 net666 vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__A2 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10115__A1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11312__A0 _06469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07531__A2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__A _04178_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14819_ clknet_leaf_32_wb_clk_i net1874 _01184_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09808__A1 _02923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\] net959 net917
+ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__a221o_1
XANTENNA__07819__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ net1230 team_03_WB.instance_to_wrap.core.register_file.registers_state\[183\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[151\] net969 net920
+ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08492__B1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[946\] net752
+ net1011 _03163_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07153_ net1190 team_03_WB.instance_to_wrap.core.register_file.registers_state\[480\]
+ net882 _03094_ net1126 vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a311o_1
XANTENNA__07047__A1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07084_ net1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[545\]
+ net895 vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08547__A1 net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A net578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_A net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06869__B team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout489_A _06779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13048__A net1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[976\]
+ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09960__S net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ _03759_ _04893_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__a21oi_1
X_06937_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[740\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[708\]
+ net769 vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout656_A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09656_ _05296_ _05597_ _05303_ _05285_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__o211a_1
XANTENNA__08576__S net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\] vssd1 vssd1 vccd1
+ vccd1 _02810_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _04545_ _04546_ _04547_ _04548_ net859 net938 vssd1 vssd1 vccd1 vccd1 _04549_
+ sky130_fd_sc_hd__mux4_1
X_09587_ net541 _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout823_A _06558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08158__S0 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08538_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[862\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[894\] net1065
+ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10200__A _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11015__B _06468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[444\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[412\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[316\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[284\]
+ net953 net1065 vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__mux4_1
XFILLER_0_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11730__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ net131 net1027 net903 net1920 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a22o_1
XANTENNA__10290__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11480_ net506 net631 _06604_ net400 net2225 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a32o_1
XANTENNA__07038__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10431_ _06020_ _06022_ _06061_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09983__A0 _05868_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ net1383 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
X_10362_ team_03_WB.instance_to_wrap.core.pc.current_pc\[22\] _06146_ vssd1 vssd1
+ vccd1 vccd1 _06195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07994__C1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ net636 _06675_ net475 net445 net1754 vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10293_ team_03_WB.instance_to_wrap.core.pc.current_pc\[5\] team_03_WB.instance_to_wrap.core.pc.current_pc\[4\]
+ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__and4_1
X_13081_ net1357 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XANTENNA__08538__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ _06773_ net482 net368 net2332 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__a22o_1
Xhold190 team_03_WB.instance_to_wrap.CPU_DAT_I\[10\] vssd1 vssd1 vccd1 vccd1 net1774
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07882__C net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11542__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__C1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10896__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout670 net674 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 _05915_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_2
Xfanout692 _02839_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
X_13983_ clknet_leaf_115_wb_clk_i _01747_ _00348_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12797__A net1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ net1411 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
XANTENNA__08486__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08171__C1 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ net1266 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
X_14604_ clknet_leaf_7_wb_clk_i _02368_ _00969_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[958\]
+ sky130_fd_sc_hd__dfstp_1
X_11816_ _06644_ net483 net330 net2185 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12796_ net1350 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14535_ clknet_leaf_66_wb_clk_i _02299_ _00900_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07277__A1 net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11747_ net648 _06569_ net456 net337 net2043 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10820__A2 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14466_ clknet_leaf_129_wb_clk_i _02230_ _00831_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _06720_ net385 net344 net2274 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13417_ net1403 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09569__A3 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08226__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ net1753 team_03_WB.instance_to_wrap.CPU_DAT_O\[0\] net837 vssd1 vssd1 vccd1
+ vccd1 _02499_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14397_ clknet_leaf_68_wb_clk_i _02161_ _00762_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09974__A0 _03488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__A1 net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13348_ net1294 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10584__B2 _02888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ net1396 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15018_ clknet_leaf_40_wb_clk_i _02738_ _01383_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09346__A _04148_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11087__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07201__A1 net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07840_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[682\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[650\]
+ net759 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12089__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14295__CLK clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ net1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[876\]
+ net888 _03710_ net1153 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__o311a_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06960__B1 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ net581 _05451_ net358 vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11836__A1 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10939__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09441_ _04826_ _05382_ net558 vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11116__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _04382_ _05312_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ net854 _04261_ _04263_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08254_ _04194_ _04195_ net855 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06871__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[1\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07205_ net1161 team_03_WB.instance_to_wrap.core.register_file.registers_state\[338\]
+ net752 team_03_WB.instance_to_wrap.core.register_file.registers_state\[370\] net1116
+ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__o221a_1
XFILLER_0_6_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12013__A1 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08217__B1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08185_ net850 _04125_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__or3_1
XFILLER_0_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout404_A _06752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1146_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08768__A1 net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07136_ net1104 team_03_WB.instance_to_wrap.core.register_file.registers_state\[960\]
+ net799 team_03_WB.instance_to_wrap.core.register_file.registers_state\[992\] net1126
+ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10575__B2 _05885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__C1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07067_ net1091 team_03_WB.instance_to_wrap.core.register_file.registers_state\[34\]
+ net894 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11001__D net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput240 net240 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput251 net251 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput262 net262 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_80_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09717__B1 _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__C1 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10878__A2 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08940__A1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07743__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ net1099 team_03_WB.instance_to_wrap.core.register_file.registers_state\[240\]
+ net897 vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout940_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08379__S0 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _04150_ _04210_ _05014_ _05071_ net559 net574 vssd1 vssd1 vccd1 vccd1 _05650_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__13662__CLK clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ team_03_WB.instance_to_wrap.core.decoder.inst\[8\] net1246 net1015 vssd1
+ vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__and3_4
X_09639_ _05356_ _05577_ _05578_ _05580_ _05575_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07223__B net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ net1257 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14018__CLK clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11601_ _06527_ net2305 net454 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12581_ net1276 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XANTENNA__10865__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ clknet_leaf_113_wb_clk_i _02084_ _00685_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13241__A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ net277 net643 net707 net698 vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and4_1
XANTENNA__10802__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire323 _05927_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
XFILLER_0_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14251_ clknet_leaf_36_wb_clk_i _02015_ _00616_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[605\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12004__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ net499 net627 _06588_ net398 net1938 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14168__CLK clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ net1422 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08759__A1 net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _06236_ _06237_ team_03_WB.instance_to_wrap.core.pc.current_pc\[13\] net678
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14182_ clknet_leaf_86_wb_clk_i _01946_ _00547_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[536\]
+ sky130_fd_sc_hd__dfrtp_1
X_11394_ net510 net637 _06749_ net407 net1996 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__a32o_1
XANTENNA__09420__A2 _02804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13133_ net1302 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
XANTENNA__07431__A1 net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ _06110_ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13064_ net1351 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10276_ _03822_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11515__A0 _06630_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07719__C1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1410 net1412 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__buf_4
X_12015_ _06763_ net480 net367 net2495 vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a22o_1
Xfanout1421 net1422 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__buf_4
Xfanout1432 net1433 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07734__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13966_ clknet_leaf_70_wb_clk_i _01730_ _00331_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10759__B _06294_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08144__C1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ net1269 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XANTENNA__11294__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08695__B1 net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ clknet_leaf_67_wb_clk_i _01661_ _00262_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09892__C1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ net1428 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ net1271 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08998__A1 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13151__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ clknet_leaf_87_wb_clk_i _02282_ _00883_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[872\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14449_ clknet_leaf_94_wb_clk_i _02213_ _00814_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12990__A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10006__A0 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold904 team_03_WB.instance_to_wrap.core.register_file.registers_state\[772\] vssd1
+ vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold915 team_03_WB.instance_to_wrap.core.register_file.registers_state\[559\] vssd1
+ vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 team_03_WB.instance_to_wrap.core.register_file.registers_state\[499\] vssd1
+ vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold937 team_03_WB.instance_to_wrap.core.register_file.registers_state\[209\] vssd1
+ vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07422__A1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\] vssd1
+ vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09990_ _05875_ net2112 net288 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold959 team_03_WB.instance_to_wrap.core.register_file.registers_state\[453\] vssd1
+ vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08941_ net1213 _04881_ _04882_ net1070 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o211a_1
XANTENNA__11506__A0 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ _04808_ _04811_ _04812_ net592 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07186__B1 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ net1078 team_03_WB.instance_to_wrap.core.register_file.registers_state\[74\]
+ net786 team_03_WB.instance_to_wrap.core.register_file.registers_state\[106\] net740
+ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07754_ net1085 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\]
+ net889 _03695_ net1143 vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__o311a_1
XANTENNA__09478__A2 _04476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07489__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[702\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\] net759 net726
+ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout354_A net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__B net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__B1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _05360_ _05365_ net555 vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__mux2_1
XANTENNA__08781__S0 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11037__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _03947_ _05148_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout521_A net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout619_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_A net1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08306_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[440\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[408\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[312\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[280\]
+ net983 net1075 vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09286_ _04922_ _05225_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__or2_1
XANTENNA__11993__A0 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__B1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08155__A team_03_WB.instance_to_wrap.core.decoder.inst\[19\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08237_ net437 net430 _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__or3b_2
XANTENNA_fanout1430_A net1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08168_ net1055 _04108_ _04109_ _04107_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout890_A net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_108_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07949__C1 net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11745__B1 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout988_A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07413__A1 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ net611 _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10624__S net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ _04037_ _04040_ net817 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12405__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _04415_ _02767_ net671 vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__mux2_1
XANTENNA__07335__A1_N net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15089__1470 vssd1 vssd1 vccd1 vccd1 _15089__1470/HI net1470 sky130_fd_sc_hd__conb_1
X_10061_ net24 net1035 net909 team_03_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1
+ vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07716__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__A1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__B1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13820_ clknet_leaf_119_wb_clk_i _01584_ _00185_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07234__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ clknet_leaf_73_wb_clk_i _01515_ _00116_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11276__A2 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ net686 _05798_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12702_ net1384 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XANTENNA__10484__B1 net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13682_ clknet_leaf_100_wb_clk_i _01446_ _00047_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08764__S net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10894_ net300 net2592 net523 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11028__A2 net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12633_ net1354 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XANTENNA__08429__B1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__A0 _05068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ net1320 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08065__A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11984__A0 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14303_ clknet_leaf_121_wb_clk_i _02067_ _00668_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[657\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ _06630_ net2803 net396 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07652__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07400__C net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12495_ net1410 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14234_ clknet_leaf_22_wb_clk_i _01998_ _00599_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11446_ net276 net643 net707 net825 vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__and4_1
XFILLER_0_81_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11736__B1 _06808_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07404__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14165_ clknet_leaf_90_wb_clk_i _01929_ _00530_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[519\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11377_ net714 net297 net698 vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13116_ net1350 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_10328_ _02767_ _06151_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14096_ clknet_leaf_81_wb_clk_i _01860_ _00461_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ net1415 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
X_10259_ _04030_ _06099_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08939__S net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08904__A1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1241 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_4
Xfanout1251 net1270 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
XANTENNA__10711__A1 _05499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__B1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1273 net1274 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_4
Xfanout1284 net1286 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_4
Xfanout1295 net1433 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_4
XANTENNA__08117__C1 net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14998_ clknet_leaf_107_wb_clk_i net46 _01363_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_13949_ clknet_leaf_60_wb_clk_i _01713_ _00314_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_92_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07470_ net1173 team_03_WB.instance_to_wrap.core.register_file.registers_state\[565\]
+ net874 vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07891__A1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _04538_ _05074_ _04779_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__or3b_4
XANTENNA__10936__C net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11975__A0 _06405_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14483__CLK clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09071_ net440 net431 _05012_ net554 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o31a_1
XANTENNA__11113__B _06541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08840__B1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ net1167 team_03_WB.instance_to_wrap.core.register_file.registers_state\[49\]
+ net873 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold701 team_03_WB.instance_to_wrap.core.register_file.registers_state\[101\] vssd1
+ vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 team_03_WB.instance_to_wrap.core.register_file.registers_state\[697\] vssd1
+ vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10952__B _05768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold723 team_03_WB.instance_to_wrap.core.register_file.registers_state\[353\] vssd1
+ vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 team_03_WB.instance_to_wrap.core.register_file.registers_state\[700\] vssd1
+ vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 team_03_WB.instance_to_wrap.core.register_file.registers_state\[231\] vssd1
+ vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 team_03_WB.instance_to_wrap.core.register_file.registers_state\[878\] vssd1
+ vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold767 team_03_WB.instance_to_wrap.core.register_file.registers_state\[147\] vssd1
+ vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07319__A net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold778 team_03_WB.instance_to_wrap.core.register_file.registers_state\[310\] vssd1
+ vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09973_ _03458_ net1837 net294 vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__mux2_1
Xhold789 team_03_WB.instance_to_wrap.core.register_file.registers_state\[457\] vssd1
+ vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11486__D net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ net1233 team_03_WB.instance_to_wrap.core.register_file.registers_state\[139\]
+ net977 team_03_WB.instance_to_wrap.core.register_file.registers_state\[171\] net938
+ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__o221a_1
XANTENNA__07159__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1011_A _02869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A _02786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[544\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[512\]
+ net986 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__mux2_1
XANTENNA__07980__C net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout471_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A _03025_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07806_ _03744_ _03747_ net814 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13056__A net1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08786_ net1054 team_03_WB.instance_to_wrap.core.register_file.registers_state\[834\]
+ net1009 team_03_WB.instance_to_wrap.core.register_file.registers_state\[866\] net1206
+ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a221o_1
XANTENNA__08108__C1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11258__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ team_03_WB.instance_to_wrap.core.decoder.inst\[13\] net1012 _03107_ vssd1
+ vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12895__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1380_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08584__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ net1164 team_03_WB.instance_to_wrap.core.register_file.registers_state\[94\]
+ net758 team_03_WB.instance_to_wrap.core.register_file.registers_state\[126\] net725
+ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__o221a_1
XANTENNA__06893__A team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09407_ net551 _04237_ _04325_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14826__CLK clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10619__S net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[473\]
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09338_ _05196_ _05202_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11966__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07634__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09269_ net588 _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__D_N _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ _06609_ net2856 net412 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12280_ net1362 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08809__S1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ _06545_ net2004 net492 vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07229__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ net703 net271 net695 vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__and3_1
XANTENNA__14206__CLK clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _05952_ _05953_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ net829 net300 vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__and2_2
XFILLER_0_101_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08347__C1 net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net12 net1035 net908 team_03_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1
+ vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
X_14921_ clknet_leaf_126_wb_clk_i _02676_ _01286_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08898__B1 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 _02632_ vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold61 team_03_WB.instance_to_wrap.core.register_file.registers_state\[980\] vssd1
+ vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 team_03_WB.instance_to_wrap.core.register_file.registers_state\[954\] vssd1
+ vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14356__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14852_ clknet_leaf_53_wb_clk_i net1790 _01217_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold83 team_03_WB.instance_to_wrap.core.register_file.registers_state\[956\] vssd1
+ vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1012\] vssd1
+ vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ clknet_leaf_46_wb_clk_i _01567_ _00168_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[157\]
+ sky130_fd_sc_hd__dfrtp_1
X_14783_ clknet_leaf_32_wb_clk_i _02547_ _01148_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10102__B _05945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _06754_ net470 net450 net2379 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11913__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13734_ clknet_leaf_75_wb_clk_i _01498_ _00099_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10946_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[5\] net308 net684 vssd1
+ vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07322__B1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13665_ clknet_leaf_2_wb_clk_i _01429_ _00030_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10877_ net273 net2210 net521 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12616_ net1351 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
X_13596_ net1274 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11957__B1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12547_ net1267 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
XANTENNA__11421__A2 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1386 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__A3 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__C_N net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12478_ net1384 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ clknet_leaf_67_wb_clk_i _01981_ _00582_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[571\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11429_ net269 net2740 net403 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15197_ net910 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_1
XANTENNA__07389__B1 _02871_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11185__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ clknet_leaf_20_wb_clk_i _01912_ _00513_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ clknet_leaf_116_wb_clk_i _01843_ _00444_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[433\]
+ sky130_fd_sc_hd__dfrtp_1
X_06970_ net1037 _02910_ _02911_ net1011 _02909_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_1392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_22 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_4
XFILLER_0_101_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
X_08640_ _04580_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1092 net1105 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ net1225 team_03_WB.instance_to_wrap.core.register_file.registers_state\[349\]
+ net961 team_03_WB.instance_to_wrap.core.register_file.registers_state\[381\] net1067
+ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07522_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[934\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[902\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[806\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\]
+ net775 net1124 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08510__C1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07864__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07453_ net1172 team_03_WB.instance_to_wrap.core.register_file.registers_state\[181\]
+ net888 net1118 vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11124__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14999__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07384_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[479\]
+ net770 team_03_WB.instance_to_wrap.core.register_file.registers_state\[511\] net1146
+ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11948__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__C _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ _05061_ _05062_ _05063_ _05064_ net856 net916 vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1059_A net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09054_ net1215 _04993_ _04994_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__and3_1
XANTENNA__11963__A3 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08005_ _03945_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or2_2
XFILLER_0_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold520 team_03_WB.instance_to_wrap.core.ru.prev_busy vssd1 vssd1 vccd1 vccd1 net2104
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold531 team_03_WB.instance_to_wrap.core.register_file.registers_state\[38\] vssd1
+ vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 team_03_WB.instance_to_wrap.core.register_file.registers_state\[57\] vssd1
+ vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__C1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold553 team_03_WB.instance_to_wrap.core.register_file.registers_state\[841\] vssd1
+ vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08041__A1 _02847_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[29\] vssd1 vssd1 vccd1
+ vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 team_03_WB.instance_to_wrap.core.register_file.registers_state\[909\] vssd1
+ vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold586 team_03_WB.instance_to_wrap.core.register_file.registers_state\[425\] vssd1
+ vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 net113 vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09956_ _05882_ net1811 net294 vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08907_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[716\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[748\] net935
+ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09264__A _03682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11479__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _03137_ _04148_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout853_A net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_03_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 net2804
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 team_03_WB.instance_to_wrap.core.register_file.registers_state\[220\] vssd1
+ vssd1 vccd1 vccd1 net2815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__B1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[32\] net986
+ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or2_1
Xhold1242 team_03_WB.instance_to_wrap.core.register_file.registers_state\[188\] vssd1
+ vssd1 vccd1 vccd1 net2826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 team_03_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 net2837
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1264 team_03_WB.instance_to_wrap.core.register_file.registers_state\[92\] vssd1
+ vssd1 vccd1 vccd1 net2848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[23\] vssd1 vssd1
+ vccd1 vccd1 net2859 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 team_03_WB.instance_to_wrap.core.register_file.registers_state\[83\] vssd1
+ vssd1 vccd1 vccd1 net2870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08769_ net847 _04693_ _04702_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11733__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__B1 net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__A net1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _06406_ _06408_ net587 vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11780_ net2505 _06613_ net332 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ net1897 net530 net525 _06357_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
XANTENNA__07855__A1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ net1395 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
X_10662_ net1135 net1585 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__or2_1
XANTENNA__09057__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12401_ net1304 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_123_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07607__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ net1403 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08804__B1 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ team_03_WB.instance_to_wrap.core.ru.prev_busy _06281_ vssd1 vssd1 vccd1 vccd1
+ _06302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15120_ net1501 vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_2
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12332_ net1299 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08280__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11954__A3 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07083__A2 _03023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ net1583 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
X_12263_ net1389 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08568__C1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ clknet_leaf_103_wb_clk_i _01766_ _00367_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[356\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11214_ net2479 net490 _06681_ net500 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XANTENNA__08032__A1 net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ net1647 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__clkbuf_1
X_11145_ net2166 net418 _06649_ net505 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
XANTENNA__07240__C1 net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08489__S net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10390__A2 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ net829 net276 vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__and2_2
XFILLER_0_21_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10027_ net1136 net100 _05903_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__mux2_1
X_14904_ clknet_leaf_48_wb_clk_i _02667_ _01269_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07543__B1 net1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A _05563_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ clknet_leaf_31_wb_clk_i net2018 _01200_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
XANTENNA__07125__C net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A2 _06699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__S0 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14766_ clknet_leaf_122_wb_clk_i _02530_ _01131_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11978_ net279 net2742 net448 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__mux2_1
XANTENNA__10767__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09113__S net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ net316 net310 net319 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[8\]
+ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or4b_1
X_13717_ clknet_leaf_89_wb_clk_i _01481_ _00082_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_14697_ clknet_leaf_42_wb_clk_i _02461_ _01062_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11642__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09048__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ clknet_leaf_82_wb_clk_i _01412_ _00013_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15068__1449 vssd1 vssd1 vccd1 vccd1 _15068__1449/HI net1449 sky130_fd_sc_hd__conb_1
XANTENNA__09599__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13579_ net1310 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XANTENNA__06980__B _02893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08271__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__A3 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08271__B2 net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11158__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08559__C1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08023__A1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ _02923_ _04565_ _04821_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__o31a_1
Xfanout307 _06397_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_4
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_4
X_09741_ _05086_ _05117_ _05119_ _05110_ net558 net572 vssd1 vssd1 vccd1 vccd1 _05683_
+ sky130_fd_sc_hd__mux4_1
X_06953_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[37\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[5\]
+ net771 vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09672_ net576 _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06884_ team_03_WB.instance_to_wrap.core.decoder.inst\[30\] team_03_WB.instance_to_wrap.core.decoder.inst\[28\]
+ team_03_WB.instance_to_wrap.core.decoder.inst\[27\] _02824_ vssd1 vssd1 vccd1 vccd1
+ _02826_ sky130_fd_sc_hd__or4_1
XANTENNA__07534__B1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08731__C1 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08623_ net847 _04564_ _04551_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_136_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10958__A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A _06550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08554_ net855 _04492_ _04495_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07505_ net1096 team_03_WB.instance_to_wrap.core.register_file.registers_state\[71\]
+ net794 team_03_WB.instance_to_wrap.core.register_file.registers_state\[103\] net749
+ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08485_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[891\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[859\]
+ net989 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
XANTENNA__11633__A2 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07436_ _03375_ _03377_ net806 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout601_A _06295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07367_ net1115 _03308_ _03307_ net1130 vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__a211o_1
XFILLER_0_91_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09106_ net1042 team_03_WB.instance_to_wrap.core.register_file.registers_state\[206\]
+ net996 team_03_WB.instance_to_wrap.core.register_file.registers_state\[238\] net916
+ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a221o_1
XANTENNA__09259__A _05012_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07298_ net814 _03239_ net719 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o21ai_1
X_09037_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[944\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[912\]
+ net981 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11149__A1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold350 team_03_WB.instance_to_wrap.core.register_file.registers_state\[301\] vssd1
+ vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13769__CLK clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 team_03_WB.instance_to_wrap.core.register_file.registers_state\[174\] vssd1
+ vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold372 net196 vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold383 net109 vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11728__S net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10632__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold394 team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\] vssd1
+ vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08610__B net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout830 _06387_ vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08970__C1 net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout841 net842 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout852 _04084_ vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07507__A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _03526_ net661 vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor2_1
XANTENNA__10109__C1 _03060_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net866 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout874 net884 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11029__A net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__clkbuf_4
X_12950_ net1343 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
Xfanout896 net901 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__buf_2
Xhold1050 team_03_WB.instance_to_wrap.core.register_file.registers_state\[223\] vssd1
+ vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07525__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\] vssd1
+ vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net638 _06710_ net479 net379 net2082 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a32o_1
Xhold1072 team_03_WB.instance_to_wrap.core.register_file.registers_state\[893\] vssd1
+ vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12881_ net1312 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
Xhold1083 team_03_WB.instance_to_wrap.core.register_file.registers_state\[146\] vssd1
+ vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1094 team_03_WB.instance_to_wrap.core.register_file.registers_state\[659\] vssd1
+ vssd1 vccd1 vccd1 net2678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13244__A net1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14620_ clknet_leaf_126_wb_clk_i _02384_ _00985_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[974\]
+ sky130_fd_sc_hd__dfstp_1
X_11832_ _06668_ net480 net330 net1995 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07242__A net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ clknet_leaf_74_wb_clk_i _02315_ _00916_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07289__C1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07828__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ _06592_ net462 net337 net2176 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XANTENNA__11624__A2 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10832__A0 net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10714_ net1787 net531 net526 _06347_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a22o_1
X_13502_ net1323 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14482_ clknet_leaf_105_wb_clk_i _02246_ _00847_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[836\]
+ sky130_fd_sc_hd__dfrtp_1
X_11694_ _06736_ net392 net344 net1918 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13433_ net1425 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
X_10645_ net1212 team_03_WB.instance_to_wrap.CPU_DAT_O\[16\] net839 vssd1 vssd1 vccd1
+ vccd1 _02483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__S net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11388__A1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14544__CLK clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ net1319 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
XANTENNA__08253__A1 net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10576_ net1873 net534 net595 _05886_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15103_ net1484 vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_2
X_12315_ net1360 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07461__C1 net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13295_ net1395 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15034_ clknet_leaf_32_wb_clk_i _02754_ _01399_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12246_ net1763 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_91_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10899__A0 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__A1 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ net1682 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12323__A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08961__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11560__B2 net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11128_ net2422 net418 _06639_ net504 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__a22o_1
XANTENNA__07417__A net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11059_ net654 net706 net267 net824 vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and4_1
XANTENNA__08713__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11863__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06975__B net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14818_ clknet_leaf_60_wb_clk_i net1863 _01183_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09808__A2 _04565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07152__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11615__A2 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14749_ clknet_leaf_120_wb_clk_i _02513_ _01114_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08270_ net937 _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__A1 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08682__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06991__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07221_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[914\] net787
+ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07152_ net1102 team_03_WB.instance_to_wrap.core.register_file.registers_state\[448\]
+ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11121__B net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07083_ net611 _03023_ _02995_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11000__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11551__B2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06869__C team_03_WB.instance_to_wrap.core.control_logic.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[848\]
+ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09724_ _04816_ _05665_ net665 vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o21a_1
X_06936_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[676\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[644\]
+ net769 vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__mux2_1
XANTENNA__08857__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09655_ _05278_ _05281_ _05300_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a21o_2
XANTENNA__14417__CLK clknet_leaf_93_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[4\] _02807_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__or3b_1
XFILLER_0_59_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1293_A net1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout649_A net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[997\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[965\]
+ net973 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _04071_ _04382_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08158__S1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08537_ net1222 team_03_WB.instance_to_wrap.core.register_file.registers_state\[990\]
+ net952 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1022\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__o221a_1
XFILLER_0_4_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout816_A _02846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__C net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ net1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[476\]
+ net951 team_03_WB.instance_to_wrap.core.register_file.registers_state\[508\] net1201
+ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__o221a_1
XANTENNA__07286__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07419_ net738 _03357_ _03358_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__o32a_1
XANTENNA__10290__B2 net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08399_ net1237 team_03_WB.instance_to_wrap.core.register_file.registers_state\[601\]
+ net990 team_03_WB.instance_to_wrap.core.register_file.registers_state\[633\] net926
+ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__o221a_1
XANTENNA__10627__S net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ team_03_WB.instance_to_wrap.core.pc.current_pc\[9\] _06137_ vssd1 vssd1 vccd1
+ vccd1 _06250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12031__A2 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10361_ net305 net304 _06188_ _06193_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10042__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07994__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ net630 _06674_ net474 net445 net2013 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ net1369 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10292_ team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] team_03_WB.instance_to_wrap.core.pc.current_pc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12031_ _06772_ net476 net367 net2550 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a22o_1
Xhold180 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[5\] vssd1 vssd1 vccd1
+ vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _02581_ vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11542__A1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07746__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__C1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 net662 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
Xfanout671 net674 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout682 _03278_ vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_4
X_15067__1448 vssd1 vssd1 vccd1 vccd1 _15067__1448/HI net1448 sky130_fd_sc_hd__conb_1
XANTENNA__12098__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13982_ clknet_leaf_58_wb_clk_i _01746_ _00347_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[336\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14097__CLK clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ net1275 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08171__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08710__A2 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12864_ net1409 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14603_ clknet_leaf_37_wb_clk_i _02367_ _00968_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[957\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11058__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ net652 _06643_ net463 net331 net2007 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a32o_1
XFILLER_0_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ net1344 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10110__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11746_ _06568_ net463 net337 net2398 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
X_14534_ clknet_leaf_78_wb_clk_i _02298_ _00899_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11677_ _06719_ net388 net347 net2396 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
X_14465_ clknet_leaf_1_wb_clk_i _02229_ _00830_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13416_ net1423 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_10628_ net1722 team_03_WB.instance_to_wrap.CPU_DAT_O\[1\] net835 vssd1 vssd1 vccd1
+ vccd1 _02500_ sky130_fd_sc_hd__mux2_1
XANTENNA__08226__A1 net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14396_ clknet_leaf_128_wb_clk_i _02160_ _00761_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[750\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12022__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11230__A0 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__B2 team_03_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13347_ net1288 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
X_10559_ net1987 net534 net595 _05869_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_84_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13278_ net1396 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ clknet_leaf_56_wb_clk_i _02737_ _01382_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12229_ net1713 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09726__B2 _04820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11533__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07832__S0 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07770_ net1169 team_03_WB.instance_to_wrap.core.register_file.registers_state\[972\]
+ net761 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1004\] net1153
+ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__o221a_1
XANTENNA__12089__A2 _06656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__S net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06960__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09440_ net553 _04712_ _04740_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _04382_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor2_1
XANTENNA__11116__B net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__C net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10020__B net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08322_ _04253_ _04254_ net862 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08253_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[722\]
+ net946 team_03_WB.instance_to_wrap.core.register_file.registers_state\[754\] net929
+ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__o221a_1
XANTENNA__07673__C1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11132__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ net806 _03142_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06857__A_N team_03_WB.instance_to_wrap.core.control_logic.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08217__A1 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08184_ net1218 team_03_WB.instance_to_wrap.core.register_file.registers_state\[211\]
+ net947 team_03_WB.instance_to_wrap.core.register_file.registers_state\[243\] net929
+ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07135_ net1112 _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10575__A2 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1139_A net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07066_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[162\] net771
+ net744 _03007_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__o211a_1
Xoutput230 net230 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XFILLER_0_112_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08441__A _04382_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput241 net241 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput252 net252 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_0_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1306_A net1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12119__A_N net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout766_A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08587__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ net1186 team_03_WB.instance_to_wrap.core.register_file.registers_state\[80\]
+ net784 team_03_WB.instance_to_wrap.core.register_file.registers_state\[112\] net735
+ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__o221a_1
XANTENNA__08379__S1 net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06919_ net809 _02859_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__and3_1
XANTENNA__11288__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ _05209_ _05211_ _05276_ net591 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ net1193 team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\]
+ net880 _02872_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout933_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09638_ net565 _05579_ net326 vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09569_ _03904_ _04235_ _04820_ net1018 net1139 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11741__S net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ net296 net2551 net455 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12580_ net1306 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XANTENNA__08456__A1 net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10865__B net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__C1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11531_ net503 net625 _06643_ net486 net1808 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__a32o_1
XANTENNA__11460__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10802__A3 net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250_ clknet_leaf_3_wb_clk_i _02014_ _00615_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[604\]
+ sky130_fd_sc_hd__dfrtp_1
X_11462_ net2784 net399 _06767_ net518 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a22o_1
XANTENNA__08208__A1 _04149_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09405__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12004__A2 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ net1315 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
XANTENNA__11212__A0 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ net285 _06141_ _06233_ net678 vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14181_ clknet_leaf_107_wb_clk_i _01945_ _00546_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[535\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ net715 net267 net697 vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10566__A2 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ net1298 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
X_10344_ _05975_ _05977_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nand2_1
XANTENNA_input62_A gpio_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13063_ net1405 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10275_ _04444_ _02768_ net671 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1400 net1404 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__buf_4
X_12014_ _06762_ net483 net367 net2267 vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1411 net1412 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__buf_4
Xfanout1422 net1426 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__buf_4
XANTENNA__07195__A1 _03136_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1433 net66 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11916__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 _06680_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ clknet_leaf_108_wb_clk_i _01729_ _00330_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11818__A2 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12916_ net1322 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08695__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ clknet_leaf_18_wb_clk_i _01660_ _00261_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[250\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09910__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ net1409 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12778_ net1256 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09121__S net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14517_ clknet_leaf_72_wb_clk_i _02281_ _00882_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11729_ net2581 _06495_ net343 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14448_ clknet_leaf_80_wb_clk_i _02212_ _00813_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11203__A0 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14379_ clknet_leaf_36_wb_clk_i _02143_ _00744_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[733\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold905 team_03_WB.instance_to_wrap.core.register_file.registers_state\[917\] vssd1
+ vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10557__A2 net535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold916 team_03_WB.instance_to_wrap.core.register_file.registers_state\[527\] vssd1
+ vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A1 net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold927 team_03_WB.instance_to_wrap.core.register_file.registers_state\[123\] vssd1
+ vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09357__A _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 team_03_WB.instance_to_wrap.core.register_file.registers_state\[136\] vssd1
+ vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold949 team_03_WB.instance_to_wrap.core.register_file.registers_state\[886\] vssd1
+ vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11098__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08940_ net1044 team_03_WB.instance_to_wrap.core.register_file.registers_state\[843\]
+ net997 team_03_WB.instance_to_wrap.core.register_file.registers_state\[875\] net1059
+ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08907__C1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08871_ _04811_ _04812_ _04808_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07186__A1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ _03761_ _03763_ net801 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__06933__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07753_ net1170 team_03_WB.instance_to_wrap.core.register_file.registers_state\[460\]
+ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__or2_1
XANTENNA__08200__S net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11127__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07684_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[542\] net758
+ net739 _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09423_ net545 _04446_ _04385_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11690__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08781__S1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout347_A _06806_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13342__A net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ _05293_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1089_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07978__C net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06882__C team_03_WB.instance_to_wrap.core.decoder.inst\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ net1234 team_03_WB.instance_to_wrap.core.register_file.registers_state\[472\]
+ net983 team_03_WB.instance_to_wrap.core.register_file.registers_state\[504\] net1205
+ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__o221a_1
XFILLER_0_111_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11442__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07646__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout514_A _06448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1256_A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09966__S net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08236_ net844 _04163_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__a21o_2
XFILLER_0_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066__1447 vssd1 vssd1 vccd1 vccd1 _15066__1447/HI net1447 sky130_fd_sc_hd__conb_1
XFILLER_0_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14605__CLK clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08167_ net1219 team_03_WB.instance_to_wrap.core.register_file.registers_state\[596\]
+ net950 team_03_WB.instance_to_wrap.core.register_file.registers_state\[628\] net915
+ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__o221a_1
XANTENNA__07486__S net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ net1245 _02808_ _02818_ net1152 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_67_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ net802 _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout883_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__C1 _06399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07049_ net611 _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10060_ net27 net1035 net909 net2875 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08374__B1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__A0 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10640__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A1 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__D1 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[2\] net309 net684 vssd1
+ vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__a21o_1
X_13750_ clknet_leaf_86_wb_clk_i _01514_ _00115_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ net1381 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XANTENNA__08049__C net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10484__B2 team_03_WB.instance_to_wrap.ADR_I\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11681__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__C1 net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10893_ _06485_ _06486_ _06484_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o21a_2
X_13681_ clknet_leaf_95_wb_clk_i _01445_ _00046_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12632_ net1365 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11433__A0 net267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12563_ net1264 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07101__A1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14302_ clknet_leaf_49_wb_clk_i _02066_ _00667_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ net265 net2700 net395 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ net1338 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14285__CLK clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11445_ net503 net625 _06572_ net397 net2039 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a32o_1
X_14233_ clknet_leaf_103_wb_clk_i _01997_ _00598_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[587\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10539__A2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__S net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14164_ clknet_leaf_95_wb_clk_i _01928_ _00529_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08081__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08601__A1 net1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11376_ net500 net627 _06740_ net405 net2563 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a32o_1
XFILLER_0_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08601__B2 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10327_ _06123_ _06125_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xnor2_1
X_13115_ net1361 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14095_ clknet_leaf_96_wb_clk_i _01859_ _00460_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[449\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09905__A _05611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ net1339 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _04030_ _06099_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11646__S net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1230 net1231 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_2
X_10189_ _03460_ _06029_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__or2_1
Xfanout1252 net1255 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1263 net1270 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1274 net1277 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_4
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_4
Xfanout1296 net1297 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_4
XFILLER_0_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14997_ clknet_leaf_125_wb_clk_i net45 _01362_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.input_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13948_ clknet_leaf_129_wb_clk_i _01712_ _00313_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[302\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10786__A net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ clknet_leaf_73_wb_clk_i _01643_ _00244_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07798__C net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10778__A2 net1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09070_ net848 _04998_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08690__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08840__A1 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08021_ net1081 net887 team_03_WB.instance_to_wrap.core.register_file.registers_state\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11727__A1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13652__CLK clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold702 team_03_WB.instance_to_wrap.core.register_file.registers_state\[492\] vssd1
+ vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold713 team_03_WB.instance_to_wrap.core.register_file.registers_state\[738\] vssd1
+ vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 team_03_WB.instance_to_wrap.core.register_file.registers_state\[823\] vssd1
+ vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_03_WB.instance_to_wrap.core.register_file.registers_state\[344\] vssd1
+ vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 team_03_WB.instance_to_wrap.core.register_file.registers_state\[774\] vssd1
+ vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold757 team_03_WB.instance_to_wrap.core.register_file.registers_state\[163\] vssd1
+ vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold768 team_03_WB.instance_to_wrap.core.register_file.registers_state\[756\] vssd1
+ vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05890_ net1895 net293 vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 team_03_WB.instance_to_wrap.core.register_file.registers_state\[377\] vssd1
+ vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08923_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[11\] net998
+ net922 _04864_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__o211a_1
XANTENNA__14008__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout297_A _06513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ _04794_ _04795_ net853 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1004_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ net809 _03745_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08785_ net864 _04720_ _04726_ net847 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14158__CLK clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _03669_ _03677_ _03660_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__o21a_1
XANTENNA__08203__S0 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08659__A1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07867__C1 net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ net738 _03605_ _03606_ _03607_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout631_A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1373_A net1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_A net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ net551 _04296_ _04121_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07598_ net1194 team_03_WB.instance_to_wrap.core.register_file.registers_state\[345\]
+ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__or2_1
XANTENNA__11415__A0 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09084__A1 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ _05208_ _05211_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__and2_1
XANTENNA__11966__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ _03727_ _05150_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11430__A3 _06756_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__A_N _05718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08219_ net1059 _04158_ _04159_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or3_1
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10635__S net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ _05073_ _05120_ _05140_ _04777_ _05127_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11718__A1 _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11230_ net268 net2552 net492 vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07398__A1 net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11161_ net2665 net420 _06658_ net518 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ _04807_ net659 _05954_ _03065_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a211oi_1
XANTENNA__07944__S net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _06622_ net2264 net423 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11974__B _06751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08347__B1 net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ net14 net1032 net906 net1983 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__o22a_1
X_14920_ clknet_leaf_124_wb_clk_i _02675_ _01285_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13247__A net1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08898__A1 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_03_WB.instance_to_wrap.core.register_file.registers_state\[984\] vssd1
+ vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_03_WB.instance_to_wrap.core.register_file.registers_state\[932\] vssd1
+ vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[31\] vssd1 vssd1 vccd1
+ vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ clknet_leaf_53_wb_clk_i net1805 _01216_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
Xhold73 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1016\] vssd1
+ vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1021\] vssd1
+ vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold95 team_03_WB.instance_to_wrap.core.register_file.registers_state\[978\] vssd1
+ vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ clknet_leaf_7_wb_clk_i _01566_ _00167_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14782_ clknet_leaf_60_wb_clk_i _02546_ _01147_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.CPU_DAT_I\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09847__B1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11994_ net298 net2858 net448 vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__mux2_1
X_13733_ clknet_leaf_108_wb_clk_i _01497_ _00098_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_10945_ team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[5\] net306 vssd1 vssd1
+ vccd1 vccd1 _06529_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ clknet_leaf_132_wb_clk_i _01428_ _00029_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08076__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ _06470_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__a21oi_4
XANTENNA__11406__A0 _06434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ net1405 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09075__A1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07411__C net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13595_ net1280 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
XANTENNA__11957__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08822__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ net1346 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
XANTENNA__08822__B2 net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12477_ net1382 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14216_ clknet_leaf_35_wb_clk_i _01980_ _00581_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[570\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11428_ net513 net265 _06756_ net403 net2068 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a32o_1
XANTENNA__08015__S net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15196_ net910 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11185__A2 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14147_ clknet_leaf_23_wb_clk_i _01911_ _00512_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[501\]
+ sky130_fd_sc_hd__dfrtp_1
X_11359_ net710 net273 net695 vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__and3_1
XANTENNA__08050__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14078_ clknet_leaf_49_wb_clk_i _01842_ _00443_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13029_ net1272 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
Xfanout1071 net1076 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_4
XANTENNA__09550__A2 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_34 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11893__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 net1088 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
Xfanout1093 net1098 vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__buf_2
X_15065__1446 vssd1 vssd1 vccd1 vccd1 _15065__1446/HI net1446 sky130_fd_sc_hd__conb_1
X_08570_ net857 _04508_ _04511_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08685__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07521_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08510__B1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07452_ net1085 net889 team_03_WB.instance_to_wrap.core.register_file.registers_state\[149\]
+ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11124__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ net1180 team_03_WB.instance_to_wrap.core.register_file.registers_state\[351\]
+ net769 team_03_WB.instance_to_wrap.core.register_file.registers_state\[383\] net1122
+ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[622\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[590\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07616__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08274__C1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10963__B _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[431\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[399\]
+ team_03_WB.instance_to_wrap.core.register_file.registers_state\[303\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[271\]
+ net989 net1074 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__mux4_1
XANTENNA__10455__S net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07092__A3 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ _03934_ _03941_ net612 _03925_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__o211a_2
XFILLER_0_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11140__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold510 team_03_WB.instance_to_wrap.core.register_file.registers_state\[242\] vssd1
+ vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08026__C1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold521 net166 vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08577__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 team_03_WB.instance_to_wrap.core.register_file.registers_state\[285\] vssd1
+ vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold543 team_03_WB.instance_to_wrap.core.register_file.registers_state\[56\] vssd1
+ vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 net201 vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07049__B _02990_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\] vssd1
+ vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_03_WB.instance_to_wrap.core.register_file.registers_state\[122\] vssd1
+ vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold587 team_03_WB.instance_to_wrap.core.register_file.registers_state\[225\] vssd1
+ vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold598 team_03_WB.instance_to_wrap.core.register_file.registers_state\[178\] vssd1
+ vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _03942_ net662 vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout581_A _02992_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout679_A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__A0 _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ net1224 team_03_WB.instance_to_wrap.core.register_file.registers_state\[588\]
+ net958 team_03_WB.instance_to_wrap.core.register_file.registers_state\[620\] net917
+ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__o221a_1
XANTENNA__11479__A3 _06603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _04816_ _05827_ net663 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__o21a_1
Xhold1210 team_03_WB.instance_to_wrap.core.register_file.registers_state\[96\] vssd1
+ vssd1 vccd1 vccd1 net2794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_03_WB.instance_to_wrap.core.register_file.registers_state\[661\] vssd1
+ vssd1 vccd1 vccd1 net2805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07065__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[714\] vssd1
+ vssd1 vccd1 vccd1 net2816 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ net568 _04650_ _04774_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a211o_1
XANTENNA__11884__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1243 team_03_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1 net2827
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10203__B _05950_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_A net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1254 team_03_WB.instance_to_wrap.core.register_file.registers_state\[670\] vssd1
+ vssd1 vccd1 vccd1 net2838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 team_03_WB.instance_to_wrap.wb.curr_state\[2\] vssd1 vssd1 vccd1 vccd1 net2849
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 team_03_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1 net2860
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 team_03_WB.instance_to_wrap.core.pc.current_pc\[3\] vssd1 vssd1 vccd1 vccd1
+ net2871 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_90_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08595__S net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ net1200 _04709_ net843 vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07719_ net1174 team_03_WB.instance_to_wrap.core.register_file.registers_state\[717\]
+ net763 team_03_WB.instance_to_wrap.core.register_file.registers_state\[749\] net739
+ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__o221a_1
XANTENNA__11636__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ net1232 team_03_WB.instance_to_wrap.core.register_file.registers_state\[456\]
+ net978 team_03_WB.instance_to_wrap.core.register_file.registers_state\[488\] net1204
+ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ team_03_WB.instance_to_wrap.core.pc.current_pc\[16\] _05812_ net601 vssd1
+ vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14943__CLK clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09057__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ team_03_WB.instance_to_wrap.core.control_logic.instruction\[0\] team_03_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ net841 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12400_ net1417 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12061__A0 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07068__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ net1423 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
X_10592_ _06301_ _06292_ team_03_WB.instance_to_wrap.READ_I net1134 vssd1 vssd1 vccd1
+ vccd1 _02533_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08804__A1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__B net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12331_ net1252 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ net1411 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__inv_2
X_15050_ net1582 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XANTENNA__08568__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14001_ clknet_leaf_94_wb_clk_i _01765_ _00366_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[355\]
+ sky130_fd_sc_hd__dfrtp_1
X_11213_ _06456_ _06478_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__nor2_1
X_12193_ net1595 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11144_ net629 _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nor2_1
XANTENNA__07240__B1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11075_ _06615_ net2266 net421 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10026_ net101 net99 net102 _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__and4_1
X_14903_ clknet_leaf_48_wb_clk_i _02666_ _01268_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.pc.current_pc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09532__A2 _04354_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A1 net1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08740__B1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14834_ clknet_leaf_55_wb_clk_i _02598_ _01199_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11890__A3 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11627__B1 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08718__S1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14765_ clknet_leaf_13_wb_clk_i _02529_ _01130_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.IO_mod.data_from_mem\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11977_ _06413_ net2757 net448 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13716_ clknet_leaf_91_wb_clk_i _01480_ _00081_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_10928_ net313 net312 net321 _02781_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a31o_1
X_14696_ clknet_leaf_53_wb_clk_i _02460_ _01061_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.ADR_I\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09048__A1 net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ clknet_leaf_99_wb_clk_i _01411_ _00012_ vssd1 vssd1 vccd1 vccd1 team_03_WB.instance_to_wrap.core.register_file.registers_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ team_03_WB.instance_to_wrap.core.decoder.inst\[10\] _06389_ _06390_ vssd1
+ vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12052__A0 _06454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08256__C1 net913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ net1313 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08534__A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12529_ net1312 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11158__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09220__A1 _03280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08023__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1560 vssd1 vssd1 vccd1 vccd1 la_data_out[115] sky130_fd_sc_hd__buf_2
XFILLER_0_2_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10905__A2 _05697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_4
Xfanout319 net320 vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__buf_2
XFILLER_0_120_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_06952_ team_03_WB.instance_to_wrap.core.register_file.registers_state\[165\] team_03_WB.instance_to_wrap.core.register_file.registers_state\[133\]
+ net771 vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__mux2_1
X_09740_ _04821_ _05679_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__o21ai_1
.ends

