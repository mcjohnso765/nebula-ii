* NGSPICE file created from team_04_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_8 abstract view
.subckt sky130_fd_sc_hd__bufinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

.subckt team_04_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__13855__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10669__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _03640_ net703 _05277_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o211a_1
X_08622_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09304__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13334__B team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _04160_ _04161_ _04162_ _04163_ net785 net806 vssd1 vssd1 vccd1 vccd1 _04164_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_46_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12830__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12665__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1071_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14032__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout427_A _07656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09134__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09105_ _04712_ _04713_ _04714_ _04715_ net794 net814 vssd1 vssd1 vccd1 vccd1 _04716_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12346__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold340 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\] vssd1 vssd1
+ vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\] vssd1 vssd1
+ vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12897__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold362 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\] vssd1 vssd1
+ vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\] vssd1 vssd1
+ vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\] vssd1 vssd1
+ vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14099__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\] vssd1 vssd1
+ vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout820 net821 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout831 net838 vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__clkbuf_8
X_09938_ net644 _03783_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or2_1
Xfanout842 net843 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__clkbuf_4
Xfanout853 net858 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_2
XANTENNA__12649__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout864 net871 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_2
Xfanout875 net883 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__clkbuf_4
Xfanout886 net889 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_4
Xfanout897 net903 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__buf_4
X_09869_ net579 net570 _05252_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__o2bb2a_1
Xhold1040 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\] vssd1 vssd1
+ vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1051 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\] vssd1 vssd1
+ vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07370_ sky130_fd_sc_hd__a21o_1
Xhold1062 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\] vssd1 vssd1
+ vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _07580_ net347 net391 net2244 vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__a22o_1
Xhold1073 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\] vssd1 vssd1
+ vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\] vssd1 vssd1
+ vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11872__A3 _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1095 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\] vssd1 vssd1
+ vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13244__B _06140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] net269 net268 vssd1 vssd1 vccd1
+ vccd1 _07310_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_29_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14550_ net1184 vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__inv_2
XANTENNA__09373__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ _06191_ _07248_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ net994 _02889_ _02891_ _07691_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10713_ _05469_ _06201_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__or2_1
X_14481_ net1273 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14356__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ _07180_ _07181_ _07179_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16220_ clknet_leaf_127_wb_clk_i _01889_ _00449_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input92_A wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ _07733_ _07854_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__o21bai_1
X_10644_ net1648 net1605 _06173_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ clknet_leaf_161_wb_clk_i _01820_ _00380_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\]
+ sky130_fd_sc_hd__dfrtp_1
X_13363_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\] team_04_WB.MEM_SIZE_REG_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__or2_1
XANTENNA__09169__B net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10575_ team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] net1094 net1053 vssd1 vssd1 vccd1
+ vccd1 _06122_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15102_ net1218 vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__inv_2
X_12314_ net2258 net499 _07601_ net440 vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__a22o_1
X_16082_ clknet_leaf_8_wb_clk_i _01751_ _00311_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_13294_ _07720_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output179_A net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ net1239 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12245_ net2215 net503 _07565_ net438 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12888__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12176_ net1979 net507 _07529_ net440 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12323__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _06215_ _06218_ net539 vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__mux2_1
X_16984_ clknet_leaf_150_wb_clk_i _02653_ _01213_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09472__X _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15935_ clknet_leaf_58_wb_clk_i _01612_ _00162_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09913__A net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11848__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ _06543_ _06545_ net537 vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_60_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10009_ _05601_ _05619_ _05600_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__a21o_1
X_15866_ clknet_leaf_96_wb_clk_i _01543_ _00093_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09124__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14817_ net1150 vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__inv_2
XANTENNA__09269__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14748_ net1125 vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_48_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14679_ net1228 vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10794__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16418_ clknet_leaf_145_wb_clk_i _02087_ _00647_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16349_ clknet_leaf_131_wb_clk_i _02018_ _00578_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10733__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12879__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13329__B team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08203__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07984_ net1079 net1028 net1024 _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _05330_ _05331_ _05332_ _05333_ net797 net803 vssd1 vssd1 vccd1 vccd1 _05334_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10969__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\]
+ net961 vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09034__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _04212_ _04213_ _04214_ _04215_ net783 net805 vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1286_A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _04143_ _04144_ _04145_ _04146_ net785 net806 vssd1 vssd1 vccd1 vccd1 _04147_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08873__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__A1 _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ _04005_ _04006_ _04007_ _04008_ net824 net733 vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12408__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10360_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05529_ vssd1
+ vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__A2 _07273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__mux2_1
X_10291_ _05535_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__nor2_1
XANTENNA__10643__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ net2334 net518 _07468_ net452 vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold170 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\] vssd1 vssd1
+ vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\] vssd1 vssd1
+ vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout650 _07520_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__clkbuf_4
Xfanout661 _03634_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__buf_6
Xfanout672 _07554_ vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09499__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09043__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13981_ _04526_ net262 net598 _03324_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a31o_1
Xfanout694 _06186_ vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
X_15720_ net1294 vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__inv_2
XANTENNA__11327__X _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ net247 net2187 net318 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09594__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08171__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15651_ net1177 vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12863_ _07563_ net327 net388 net1946 vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a22o_1
XANTENNA__13047__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14602_ net1286 vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__inv_2
X_11814_ net651 net241 vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__and2_1
X_15582_ net1216 vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__inv_2
X_12794_ net220 net2443 net324 vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17321_ net1377 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_164_Left_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ net1173 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_174_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _07217_ _07218_ _07232_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_174_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09671__A1 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11503__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ net1312 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XFILLER_0_166_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_851 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14464_ net1263 vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__inv_2
XANTENNA_input95_X net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11676_ net464 _07154_ _07164_ net287 vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_12_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16203_ clknet_leaf_23_wb_clk_i _01872_ _00432_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\]
+ sky130_fd_sc_hd__dfrtp_1
X_13415_ net1084 team_04_WB.MEM_SIZE_REG_REG\[21\] vssd1 vssd1 vccd1 vccd1 _07841_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_126_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10627_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\]
+ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__or4_1
X_17183_ clknet_leaf_87_wb_clk_i _02795_ _01412_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14395_ net1255 vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14814__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16134_ clknet_leaf_19_wb_clk_i _01803_ _00363_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_13346_ _07770_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10558_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[14\]
+ _06110_ net1047 vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07985__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12554__C_N net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ clknet_leaf_141_wb_clk_i _01734_ _00294_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ _05613_ _05614_ net624 vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__o21a_1
X_10489_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] net1006 _06053_ _06063_
+ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a22o_1
XANTENNA__10780__C net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_173_Left_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15016_ net1118 vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__inv_2
XANTENNA__09119__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ net211 net673 vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_121_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12053__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12730__A1 _07455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09914__Y _05525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12159_ _05279_ _06181_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nor2_8
XFILLER_0_75_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16967_ clknet_leaf_168_wb_clk_i _02636_ _01196_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10789__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15918_ clknet_leaf_79_wb_clk_i _01595_ _00145_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16898_ clknet_leaf_146_wb_clk_i _02567_ _01127_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11288__A2_N net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15849_ clknet_leaf_94_wb_clk_i _01526_ _00076_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13038__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09789__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11049__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08693__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09370_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\]
+ net945 vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08321_ net778 _03931_ net762 vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ net643 _03861_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12228__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12549__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08183_ _03790_ _03791_ _03792_ _03793_ net832 net737 vssd1 vssd1 vccd1 vccd1 _03794_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12943__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_160_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_171_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11757__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11221__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08281__X _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11772__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09029__S net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_15__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10732__A0 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08868__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout661_A _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10699__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _05313_ _05314_ _05315_ _05316_ net797 net803 vssd1 vssd1 vccd1 vccd1 _05317_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12485__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] vssd1
+ vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09637_ net719 _05247_ _05236_ _05235_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13029__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_A _03555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ net731 _05172_ net714 vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08519_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\]
+ net846 vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10638__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09653__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ net767 _05109_ _05098_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ net569 _06217_ _06272_ net365 _05031_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__o32a_1
XFILLER_0_37_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08861__C1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11461_ net630 _04865_ net358 vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13200_ _03548_ _07687_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__nand2_4
X_10412_ _05734_ _05739_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__xor2_1
X_14180_ _03393_ _03394_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[5\]
+ sky130_fd_sc_hd__nor2_1
X_11392_ _06863_ _06880_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09728__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13131_ _07565_ net369 net294 net1933 vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10343_ _05531_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input55_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ net2656 net1055 _05869_ _05872_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__a22o_1
X_13062_ _07283_ net2445 net303 vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__mux2_1
XANTENNA__11993__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ net236 net680 vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_167_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08778__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16821_ clknet_leaf_12_wb_clk_i _02490_ _01050_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout480 net494 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 net494 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
X_16752_ clknet_leaf_190_wb_clk_i _02421_ _00981_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\]
+ sky130_fd_sc_hd__dfrtp_1
X_13964_ net152 net1064 vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__and2_1
X_15703_ net1258 vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__inv_2
X_12915_ _07617_ net342 net386 net2063 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a22o_1
X_16683_ clknet_leaf_31_wb_clk_i _02352_ _00912_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\]
+ sky130_fd_sc_hd__dfrtp_1
X_13895_ _03169_ _03195_ _03269_ _03243_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09828__A_N _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15634_ net1176 vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ _07544_ net330 net392 net1956 vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a22o_1
XANTENNA__14312__S1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09402__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__A1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15565_ net1144 vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__inv_2
X_12777_ _07504_ net338 net396 net1869 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a22o_1
XANTENNA__12329__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17304_ net1360 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XFILLER_0_150_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11233__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14516_ net1192 vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11728_ _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__or2_1
XANTENNA__11451__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15496_ net1117 vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ net1401 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
X_14447_ net1276 vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _06530_ _06949_ _06886_ _06537_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a2bb2o_1
X_17166_ clknet_leaf_93_wb_clk_i _02778_ _01395_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_14378_ net1453 vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07958__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold906 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\] vssd1 vssd1
+ vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\] vssd1 vssd1
+ vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ clknet_leaf_33_wb_clk_i _01786_ _00346_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\]
+ sky130_fd_sc_hd__dfrtp_1
X_13329_ net1086 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 _07755_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_24_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold928 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\] vssd1 vssd1
+ vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
X_17097_ clknet_leaf_91_wb_clk_i _02732_ _01326_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold939 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\] vssd1 vssd1
+ vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16048_ clknet_leaf_0_wb_clk_i _01717_ _00277_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12351__X _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13607__B _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12938__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10493__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout242_A _07295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08304_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__mux2_1
XANTENNA__11143__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09284_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__mux2_1
XANTENNA__12673__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13996__C _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11797__B _07280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\]
+ net946 vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08452__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08097_ _03704_ _03705_ _03706_ _03707_ net785 net800 vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload90 clknet_leaf_144_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09246__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11902__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09283__A net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08999_ net768 _04609_ _04598_ _04597_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__o2bb2a_4
Xclkbuf_leaf_188_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_188_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10961_ _06364_ _06367_ _06449_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net2254 net404 net327 _07302_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a22o_1
XANTENNA__09730__B _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _07116_ net274 _06175_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__o21ai_1
X_10892_ _04947_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__nor2_1
XANTENNA__09222__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ _07602_ net479 net408 net2060 vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ net1222 vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__inv_2
XANTENNA__12630__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12562_ _07529_ net481 net416 net1727 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13973__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ _03463_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11513_ net632 net630 net628 net627 net546 net539 vssd1 vssd1 vccd1 vccd1 _07002_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11988__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15281_ net1270 vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__inv_2
XANTENNA__10892__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ _07490_ net483 net425 net2128 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13186__A1 _07622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17020_ clknet_leaf_127_wb_clk_i _02689_ _01249_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\]
+ sky130_fd_sc_hd__dfrtp_1
X_14232_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] _03422_ vssd1
+ vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11444_ team_04_WB.MEM_SIZE_REG_REG\[16\] _06508_ vssd1 vssd1 vccd1 vccd1 _06933_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09485__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08288__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] _03368_
+ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_169_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11375_ _06427_ _06444_ _06448_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ _07546_ net379 net300 net1758 vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a22o_1
X_10326_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\] _05531_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21oi_1
X_14094_ net1458 _06134_ net1034 vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ _07506_ net370 net306 net1647 vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a22o_1
X_10257_ _05537_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__or2_1
XANTENNA__12697__B1 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1220 net1254 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
Xfanout1231 net1234 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_4
X_10188_ net622 _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor2_1
XANTENNA__08301__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_2
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
Xfanout1264 net1297 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__buf_4
XANTENNA__10172__B2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12331__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1275 net1279 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__clkbuf_4
X_16804_ clknet_leaf_173_wb_clk_i _02473_ _01033_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_14__f_wb_clk_i_X clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1286 net1288 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_4
Xfanout1297 net35 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_4
X_14996_ net1214 vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__inv_2
XANTENNA__08117__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13947_ net160 net1064 vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__and2_1
X_16735_ clknet_leaf_156_wb_clk_i _02404_ _00964_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\]
+ sky130_fd_sc_hd__dfrtp_1
X_16666_ clknet_leaf_38_wb_clk_i _02335_ _00895_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\]
+ sky130_fd_sc_hd__dfrtp_1
X_13878_ _02932_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__and2_1
XANTENNA__08537__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09132__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07971__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15617_ net1131 vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__inv_2
X_12829_ _07527_ net333 net393 net1595 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a22o_1
X_16597_ clknet_leaf_15_wb_clk_i _02266_ _00826_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12059__A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15548_ net1145 vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__inv_2
XANTENNA__08971__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12621__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11898__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15479_ net1230 vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08020_ _03607_ _03630_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nor2_4
XFILLER_0_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17218_ net1424 _02828_ _01463_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold703 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\] vssd1 vssd1
+ vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ clknet_leaf_85_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[3\]
+ _01378_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_141_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold714 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\] vssd1 vssd1
+ vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold725 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\] vssd1 vssd1
+ vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\] vssd1 vssd1
+ vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14126__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold747 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\] vssd1 vssd1
+ vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold758 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\] vssd1 vssd1
+ vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net635 _04612_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold769 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\] vssd1 vssd1
+ vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08922_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08853_ net726 _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08451__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08784_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\]
+ net866 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_140_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12668__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10977__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10696__B net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09042__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ net731 _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09608__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ net767 _04946_ _04935_ _04929_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_146_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12612__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13955__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__A1 _07604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__mux2_1
X_09198_ _04805_ _04806_ _04807_ _04808_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04809_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08149_ _03756_ _03757_ _03758_ _03759_ net786 net807 vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_75_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14912__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08595__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11160_ _03920_ net363 _06648_ net582 vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] _05058_ vssd1
+ vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_8_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11091_ net627 net547 _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__a21o_1
XANTENNA__12432__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_164_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _05551_ _05652_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or2_1
XANTENNA__09217__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08442__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold52 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\] vssd1 vssd1
+ vccd1 vccd1 net1489 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ net1217 vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__inv_2
Xhold63 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold74 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\] vssd1 vssd1 vccd1
+ vccd1 net1511 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 _02762_ vssd1 vssd1 vccd1 vccd1 net1522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13801_ _03190_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__or2_1
Xhold96 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[19\] vssd1 vssd1
+ vccd1 vccd1 net1533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A DAT_I[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ net1154 vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
XANTENNA__10887__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ net211 net681 vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__and2_1
XANTENNA__14359__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ clknet_leaf_113_wb_clk_i _02189_ _00749_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\]
+ sky130_fd_sc_hd__dfrtp_1
X_13732_ _06992_ net271 net710 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10944_ _04865_ _06428_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__xnor2_2
XANTENNA__12851__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16451_ clknet_leaf_118_wb_clk_i _02120_ _00680_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13663_ team_04_WB.ADDR_START_VAL_REG\[3\] _03046_ _03053_ vssd1 vssd1 vccd1 vccd1
+ _03054_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10875_ _06362_ _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__nor2_1
X_15402_ net1105 vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ _07583_ net490 net414 net2178 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
XANTENNA__11406__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08791__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16382_ clknet_leaf_158_wb_clk_i _02051_ _00611_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12603__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ net1093 _02984_ net1045 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_54_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_85_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ net1110 vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08283__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12545_ net2441 net249 net423 vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13915__A1_N _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15264_ net1210 vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12476_ net608 net224 net683 vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__and3_1
XANTENNA__08092__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17003_ clknet_leaf_17_wb_clk_i _02672_ _01232_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\]
+ sky130_fd_sc_hd__dfrtp_1
X_14215_ _03416_ _03364_ _03415_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[6\]
+ sky130_fd_sc_hd__and3b_1
X_11427_ team_04_WB.MEM_SIZE_REG_REG\[11\] team_04_WB.MEM_SIZE_REG_REG\[10\] _06504_
+ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__and3_1
XANTENNA__08035__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15195_ net1136 vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14108__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _03365_ _03367_ _03360_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[0\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ net571 _06609_ _06846_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__o21ba_1
XANTENNA__10393__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08050__A3 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08681__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _05533_ vssd1
+ vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__xor2_2
XANTENNA__10561__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ net1473 _06100_ net1032 vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__mux2_1
X_11289_ _04477_ net363 _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_5_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13028_ _07489_ net369 net306 net2301 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a22o_1
XANTENNA__09630__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1050 _06075_ vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__buf_2
Xfanout1061 _03351_ vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__buf_2
Xfanout1072 net1073 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11893__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_2
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__buf_2
XFILLER_0_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13095__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__A _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ net1165 vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16718_ clknet_leaf_30_wb_clk_i _02387_ _00947_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12842__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16649_ clknet_leaf_123_wb_clk_i _02318_ _00878_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09121_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__mux2_1
XANTENNA__13620__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12076__X _07493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08206__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12236__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ _03599_ _03604_ _03608_ _03612_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or4b_1
Xhold500 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\] vssd1 vssd1
+ vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12951__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold511 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\] vssd1 vssd1
+ vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold522 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\] vssd1 vssd1
+ vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\] vssd1 vssd1
+ vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\] vssd1 vssd1
+ vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 net112 vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold566 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\] vssd1 vssd1
+ vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\] vssd1 vssd1
+ vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13348__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold588 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\] vssd1 vssd1
+ vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09954_ net638 _04275_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold599 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\] vssd1 vssd1
+ vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1114_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09037__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__mux2_1
XANTENNA__08800__A1_N net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _04440_ _04474_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__nor2_1
Xhold1200 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\] vssd1 vssd1
+ vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\] vssd1
+ vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1222 net164 vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ _03503_ net1008 net1007 _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a32o_1
XANTENNA__10687__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08876__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08767_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12833__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__mux2_1
XANTENNA__08501__A1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10660_ net2662 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1
+ vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09500__S net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11939__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09319_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__mux2_1
X_10591_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[3\]
+ _06132_ net1049 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12061__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ net2059 net502 _07609_ net459 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a22o_1
XANTENNA__08360__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08116__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15738__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ net2393 net505 _07573_ net451 vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
XANTENNA__13010__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14642__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14000_ _05445_ _03308_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nor2_1
XANTENNA__09765__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ net288 _06693_ _06697_ _06700_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12192_ net2284 net508 _07537_ net446 vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10375__B2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11143_ net555 _06213_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_132_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15951_ clknet_leaf_86_wb_clk_i net1804 _00178_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.prev_BUSY_O
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09174__C _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ net665 _05375_ _05340_ _03781_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a211o_1
XANTENNA__08415__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11324__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _05579_ _05581_ _05634_ _05580_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__a31o_1
X_14902_ net1224 vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__inv_2
X_15882_ clknet_leaf_73_wb_clk_i _01559_ _00109_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13077__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ net1270 vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14764_ net1128 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__inv_2
X_11976_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] net760 _03631_
+ _07434_ net696 vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__a221o_1
XANTENNA__12824__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ net1001 _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16503_ clknet_leaf_167_wb_clk_i _02172_ _00732_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ net579 _06402_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14695_ net1143 vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13646_ _07130_ _07216_ _07687_ _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__a22o_1
X_16434_ clknet_leaf_9_wb_clk_i _02103_ _00663_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ _04246_ _06299_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09410__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16365_ clknet_leaf_40_wb_clk_i _02034_ _00594_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13577_ _02965_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__nor2_1
XANTENNA__10556__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12052__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12337__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10789_ net587 _06250_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_54_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11241__A team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15316_ net1225 vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12528_ net2386 net226 net420 vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16296_ clknet_leaf_118_wb_clk_i _01965_ _00525_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15247_ net1196 vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13001__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ net2431 net428 _07649_ net519 vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08103__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ net1111 vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11563__B1 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14129_ team_04_WB.MEM_SIZE_REG_REG\[28\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[28\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__o221a_1
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12072__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 _07680_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12107__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13455__X _02846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_77_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10669__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _03637_ _05279_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08621_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
XANTENNA__13068__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908__1 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__inv_2
XFILLER_0_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__mux2_1
XANTENNA__12815__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17319__1375 vssd1 vssd1 vccd1 vccd1 _17319__1375/HI net1375 sky130_fd_sc_hd__conb_1
XFILLER_0_166_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08483_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__mux2_1
XANTENNA__12946__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07900__Y _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13240__A0 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout322_A _07671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1064_A net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09104_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12594__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__mux2_1
XANTENNA__12681__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13543__A1 _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09556__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12346__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold330 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\] vssd1 vssd1
+ vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\] vssd1 vssd1
+ vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout789_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\] vssd1 vssd1
+ vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold374 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\] vssd1 vssd1
+ vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\] vssd1 vssd1
+ vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\] vssd1 vssd1
+ vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 net811 vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
Xfanout821 _03419_ vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_2
X_09937_ _05546_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__nor2_1
Xfanout832 net838 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net859 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout956_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout854 net855 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__clkbuf_4
Xfanout865 net871 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11857__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout876 net883 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__clkbuf_4
Xfanout887 net889 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
X_09868_ net625 net556 vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__nand2_1
Xhold1030 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\] vssd1 vssd1
+ vccd1 vccd1 net2467 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__clkbuf_4
XANTENNA_hold367_A team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1041 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\] vssd1 vssd1
+ vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\] vssd1 vssd1
+ vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
Xhold1063 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\] vssd1 vssd1
+ vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1074 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\] vssd1 vssd1
+ vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\]
+ net895 vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__mux2_1
Xhold1085 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\] vssd1 vssd1
+ vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11326__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ net758 _05854_ net697 _04274_ net693 vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__a221o_1
Xhold1096 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\] vssd1 vssd1
+ vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12806__A0 _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_159_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout911_X net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ _06191_ _07248_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13500_ _03496_ _05815_ net1099 vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__mux2_1
XANTENNA__11613__X _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10712_ _05442_ _05447_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14480_ net1279 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__inv_2
X_11692_ _06340_ _06343_ _06658_ net463 vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09230__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13431_ team_04_WB.MEM_SIZE_REG_REG\[26\] _07730_ _07856_ vssd1 vssd1 vccd1 vccd1
+ _07857_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13231__A0 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10643_ net1555 team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__mux2_1
XANTENNA__12034__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ clknet_leaf_14_wb_clk_i _01819_ _00379_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input85_A wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ _07786_ _07787_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_172_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10574_ _06121_ net1588 net1021 vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XANTENNA__09169__C _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15101_ net1154 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__inv_2
X_12313_ net247 net668 vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ clknet_leaf_180_wb_clk_i _01750_ _00310_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_86_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13293_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] vssd1 vssd1 vccd1
+ vccd1 _07722_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15032_ net1208 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12244_ net239 net672 vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_111_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12175_ net242 net647 vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__and2_1
X_11126_ _06612_ _06614_ net563 vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__mux2_1
X_16983_ clknet_leaf_173_wb_clk_i _02652_ _01212_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\]
+ sky130_fd_sc_hd__dfrtp_1
X_15934_ clknet_leaf_58_wb_clk_i _01611_ _00161_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfrtp_1
X_11057_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10008_ _05604_ _05618_ _05603_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_95_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15865_ clknet_leaf_96_wb_clk_i _01542_ _00092_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__07921__C1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10778__C net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14816_ net1154 vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__inv_2
XANTENNA__07978__A1_N net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14747_ net1126 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__inv_2
X_11959_ net653 net231 vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__and2_1
XANTENNA__14547__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14678_ net1223 vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09140__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13629_ _07799_ _03019_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__or2_1
X_16417_ clknet_leaf_130_wb_clk_i _02086_ _00646_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_150_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12576__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16348_ clknet_leaf_128_wb_clk_i _02017_ _00577_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16279_ clknet_leaf_161_wb_clk_i _01948_ _00508_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12328__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13525__B2 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07983_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[1\] team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nand2_1
X_09722_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__mux2_1
XANTENNA__11839__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__X _06140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09315__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ net781 _05263_ net764 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_87_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout272_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09584_ _05031_ _05086_ _05142_ _05194_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_26_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08535_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12676__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13361__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1279_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08466_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12016__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout325_X net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12567__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__C net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09018_ _04617_ _04623_ _04628_ net732 net715 vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o221a_1
X_10290_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05534_ vssd1
+ vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold160 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\] vssd1 vssd1
+ vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\] vssd1 vssd1
+ vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\] vssd1 vssd1
+ vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\] vssd1 vssd1
+ vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 net641 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_4
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_4
X_13980_ net143 net1064 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__and2_1
Xfanout673 _07554_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__buf_2
XANTENNA__09043__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 net685 vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__buf_4
Xfanout695 _06186_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_4
X_12931_ net239 net2238 net318 vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ net1177 vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__inv_2
X_12862_ _07562_ net333 net389 net2129 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14601_ net1282 vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__inv_2
X_11813_ net693 _06839_ _07294_ net615 vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__a211oi_4
X_15581_ net1154 vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
X_12793_ net214 net2304 net324 vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ net1376 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
X_14532_ net1175 vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_174_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _06627_ _06655_ _07199_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_174_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08365__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09671__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17251_ net1311 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
X_14463_ net1285 vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__inv_2
XANTENNA__11503__B _06991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11675_ _06280_ _06967_ _07156_ _07161_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_12_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _07830_ _07833_ _07835_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__o31a_1
XFILLER_0_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12558__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16202_ clknet_leaf_164_wb_clk_i _01871_ _00431_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__or4_1
X_17182_ clknet_leaf_89_wb_clk_i _02794_ _01411_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_14394_ net1476 vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output191_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__B _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16133_ clknet_leaf_4_wb_clk_i _01802_ _00362_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] team_04_WB.MEM_SIZE_REG_REG\[9\]
+ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10557_ team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06110_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07985__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16064_ clknet_leaf_140_wb_clk_i _01733_ _00293_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_13276_ net69 net2646 net978 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08304__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17318__1374 vssd1 vssd1 vccd1 vccd1 _17318__1374/HI net1374 sky130_fd_sc_hd__conb_1
X_10488_ _06020_ _06046_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__or2_1
XANTENNA__11518__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15015_ net1134 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__inv_2
X_12227_ net701 _06194_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__or3_1
XANTENNA__09726__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12730__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ _07445_ net2590 net514 vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__mux2_1
XANTENNA__10741__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1053 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11109_ _06267_ _06596_ _06597_ net357 _03864_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__o32a_1
X_16966_ clknet_leaf_20_wb_clk_i _02635_ _01195_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\]
+ sky130_fd_sc_hd__dfrtp_1
X_12089_ net2426 net355 _07499_ net461 vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09135__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15917_ clknet_leaf_79_wb_clk_i _01594_ _00144_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16897_ clknet_leaf_134_wb_clk_i _02566_ _01126_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08793__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15848_ clknet_leaf_86_wb_clk_i _01525_ _00075_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15779_ net1287 vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08320_ _03927_ _03928_ _03929_ _03930_ net787 net801 vssd1 vssd1 vccd1 vccd1 _03931_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11454__C1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08251_ _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13746__B2 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08182_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\]
+ net883 vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11221__A2 _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput210 net210 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08214__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12244__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12721__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A3 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10732__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13356__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07966_ net772 _03567_ net762 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12260__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10699__B net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09705_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\]
+ net970 vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__mux2_1
XANTENNA__08689__A0 _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1 _03512_
+ sky130_fd_sc_hd__inv_2
XANTENNA__09886__C1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_80 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout654_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _05241_ _05246_ net724 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08884__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09567_ net724 _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout442_X net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout919_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12788__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09498_ _05103_ _05108_ net774 vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08449_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13737__B2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ _05464_ _06884_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10411_ net617 _05992_ _05616_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or3b_1
X_11391_ net753 _06879_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09728__B net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ _07564_ net371 net294 net2269 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a22o_1
X_10342_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _05530_ vssd1
+ vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__nor2_1
XANTENNA__12960__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08124__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ net218 net2521 net302 vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__mux2_1
X_10273_ net278 _05871_ net1074 vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08916__A1 _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ net2501 net515 _07459_ net443 vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XANTENNA__11993__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12712__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input48_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08392__A2 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ clknet_leaf_1_wb_clk_i _02489_ _01049_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__clkbuf_4
Xfanout481 net494 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16751_ clknet_leaf_190_wb_clk_i _02420_ _00980_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout492 net493 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_4
X_13963_ _04028_ net262 net598 _03315_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__a31o_1
XANTENNA__13673__B1 _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15702_ net1261 vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__inv_2
X_12914_ _07616_ net343 net386 net2036 vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__a22o_1
XANTENNA__11684__C1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13894_ net1592 net1067 net1042 _03272_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a22o_1
X_16682_ clknet_leaf_162_wb_clk_i _02351_ _00911_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15633_ net1174 vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _07543_ net330 net392 net1797 vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output204_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12779__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ _07503_ net346 net399 net1761 vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a22o_1
X_15564_ net1120 vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12329__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17303_ net1359 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_14_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14515_ net1192 vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__inv_2
X_11727_ net273 vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15495_ net1141 vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__inv_2
XANTENNA__11451__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ net1299 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
X_14446_ net1291 vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__inv_2
X_11658_ _04644_ net365 _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10609_ net49 net48 net51 net50 vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__or4_1
X_17165_ clknet_leaf_93_wb_clk_i _02777_ _01394_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10564__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14377_ net1455 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09638__B _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12345__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ _06407_ _06413_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold907 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\] vssd1 vssd1
+ vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
X_13328_ _07749_ _07752_ _07753_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__o21bai_1
Xhold918 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\] vssd1 vssd1
+ vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ clknet_leaf_2_wb_clk_i _01785_ _00345_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_17096_ clknet_leaf_105_wb_clk_i _02731_ _01325_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold929 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\] vssd1 vssd1
+ vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13259_ net77 team_04_WB.ADDR_START_VAL_REG\[17\] net978 vssd1 vssd1 vccd1 vccd1
+ _01647_ sky130_fd_sc_hd__mux2_1
X_16047_ clknet_leaf_186_wb_clk_i _01716_ _00276_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_23_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12703__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_73 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12467__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16949_ clknet_leaf_35_wb_clk_i _02618_ _01178_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09421_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09352_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\]
+ net893 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__mux2_1
XANTENNA__13967__A1 _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08209__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08303_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__mux2_1
X_09283_ net661 _03724_ _03835_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__and3_1
XANTENNA__12954__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14735__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10650__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08165_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\]
+ net946 vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout402_A _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1144_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08096_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13785__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload80 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__bufinv_8
XFILLER_0_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload91 clknet_leaf_145_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_101_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12155__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08879__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _04603_ _04608_ net776 vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07949_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__mux2_1
XANTENNA__13655__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_170_Right_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15805__24 clknet_leaf_42_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10960_ _06370_ _06376_ _06377_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__mux2_1
X_10891_ _04973_ _06292_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17317__1373 vssd1 vssd1 vccd1 vccd1 _17317__1373/HI net1373 sky130_fd_sc_hd__conb_1
XFILLER_0_168_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _07601_ net481 net408 net2224 vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a22o_1
XANTENNA_input102_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_157_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_157_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08119__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _07528_ net480 net416 net1857 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14300_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ _03462_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\] vssd1 vssd1
+ vccd1 vccd1 _03466_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11512_ _06206_ _06998_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__or3_1
X_15280_ net1162 vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12492_ _07489_ net485 net425 net1864 vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] _03422_ vssd1
+ vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11443_ net753 _06920_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__and3_2
XFILLER_0_124_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13186__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09485__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ _03374_ _03380_ _03379_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a21oi_1
X_11374_ _06508_ _06862_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_169_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14135__A1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ _07545_ net381 net301 net1939 vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a22o_1
X_10325_ net619 _05917_ _05915_ net282 vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a211o_1
XANTENNA__15476__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14093_ net1460 _06132_ net1034 vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__mux2_1
XANTENNA__08789__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12146__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ _07505_ net369 net306 net1649 vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a22o_1
XANTENNA__09474__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _05536_ vssd1
+ vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__nor2_1
XANTENNA__13894__B1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
Xfanout1221 net1224 vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_4
Xfanout1232 net1234 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__buf_2
X_10187_ _05669_ _05772_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__xor2_1
Xfanout1243 net1253 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_2
Xfanout1254 net35 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_4
X_16803_ clknet_leaf_123_wb_clk_i _02472_ _01032_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1265 net1280 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__buf_4
Xfanout1276 net1278 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__buf_4
Xfanout1287 net1288 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_4
XANTENNA__12449__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__A1_N net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14995_ net1227 vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11657__C1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16734_ clknet_leaf_142_wb_clk_i _02403_ _00963_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\]
+ sky130_fd_sc_hd__dfrtp_1
X_13946_ _03079_ _03305_ net103 net1071 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09413__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10559__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16665_ clknet_leaf_177_wb_clk_i _02334_ _00894_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\]
+ sky130_fd_sc_hd__dfrtp_1
X_13877_ _02930_ _02941_ _03258_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or3_1
XANTENNA__07971__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15616_ net1212 vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__inv_2
X_12828_ _07526_ net333 net393 net1594 vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a22o_1
X_16596_ clknet_leaf_3_wb_clk_i _02265_ _00825_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12059__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15547_ net1138 vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12759_ _07486_ net331 net398 net1814 vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11898__B _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15478_ net1223 vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17217_ net1423 _02827_ _01461_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14429_ net1272 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17148_ clknet_leaf_85_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[2\]
+ _01377_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold704 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\] vssd1 vssd1
+ vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\] vssd1 vssd1
+ vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\] vssd1 vssd1
+ vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold737 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\] vssd1 vssd1
+ vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ net635 _04612_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__or2_1
Xhold748 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\] vssd1 vssd1
+ vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ clknet_leaf_45_wb_clk_i _00027_ _01308_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12137__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold759 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\] vssd1 vssd1
+ vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08699__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ _03866_ _04088_ _04303_ _04531_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__nand4_4
XFILLER_0_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13885__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08852_ _04459_ _04460_ _04461_ _04462_ net836 net739 vssd1 vssd1 vccd1 vccd1 _04463_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08783_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\]
+ net866 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__mux2_1
XANTENNA__13637__B1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout352_A net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ _05011_ _05012_ _05013_ _05014_ net833 net738 vssd1 vssd1 vccd1 vccd1 _05015_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _04940_ _04945_ net777 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12684__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1261_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__mux2_1
XANTENNA__11820__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__mux2_1
XANTENNA__13168__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__B _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09197_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12376__A0 _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_X net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08044__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\]
+ net924 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__mux2_1
XANTENNA__09241__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__A1 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__B2 team_04_WB.ADDR_START_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08079_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
XANTENNA__12128__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10110_ _03500_ _05058_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08402__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ net589 net551 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__and2_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12432__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11329__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _05552_ _05651_ _05553_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__o21a_1
Xhold20 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\] vssd1 vssd1
+ vccd1 vccd1 net1457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\] vssd1 vssd1
+ vccd1 vccd1 net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\] vssd1 vssd1
+ vccd1 vccd1 net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\] vssd1 vssd1
+ vccd1 vccd1 net1501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 net140 vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ team_04_WB.ADDR_START_VAL_REG\[16\] _03189_ vssd1 vssd1 vccd1 vccd1 _03191_
+ sky130_fd_sc_hd__nor2_1
Xhold86 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[29\] vssd1 vssd1
+ vccd1 vccd1 net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1534 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ net1125 vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__inv_2
X_11992_ net701 _06194_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__or3_4
XANTENNA__08638__A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _03107_ _03109_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__or3_1
X_10943_ net632 _06430_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11335__Y _06824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12851__A1 _07549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16450_ clknet_leaf_144_wb_clk_i _02119_ _00679_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\]
+ sky130_fd_sc_hd__dfrtp_1
X_13662_ net1000 _03052_ _03049_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21oi_1
X_10874_ _06360_ _06361_ _04556_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15401_ net1134 vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__inv_2
XANTENNA__09155__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12613_ _07582_ net490 net414 net2032 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a22o_1
X_13593_ _07768_ _07815_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16381_ clknet_leaf_131_wb_clk_i _02050_ _00610_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12544_ net2315 net251 net420 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__mux2_1
XANTENNA__08902__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ net1169 vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08283__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13159__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12475_ net2533 net430 _07650_ net524 vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
X_15263_ net1249 vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__inv_2
XANTENNA__12367__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input70_X net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17002_ clknet_leaf_166_wb_clk_i _02671_ _01231_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\]
+ sky130_fd_sc_hd__dfrtp_1
X_14214_ _03521_ _03413_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__nor2_1
XANTENNA__08035__A1 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ net462 _06905_ _06909_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__o22a_2
XFILLER_0_34_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12906__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15194_ net1137 vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _03522_ _03366_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ net567 _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ _05900_ _05902_ net279 vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09408__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ net1465 _06098_ net1034 vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__mux2_1
XANTENNA__17194__Q team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11288_ _04476_ net362 net357 _04475_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13867__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ _07488_ net377 net308 net1870 vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a22o_1
XANTENNA__11239__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ _05683_ _05764_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1040 net1042 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09630__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1051 net1054 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__buf_2
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1062 _03350_ vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__buf_2
Xfanout1073 _07700_ vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__clkbuf_4
Xfanout1084 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 net1084 sky130_fd_sc_hd__clkbuf_2
Xfanout1095 net1097 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__buf_2
XFILLER_0_156_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14978_ net1240 vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__inv_2
X_16717_ clknet_leaf_32_wb_clk_i _02386_ _00946_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\]
+ sky130_fd_sc_hd__dfrtp_1
X_13929_ _03015_ _03094_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15796__15 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__inv_2
XFILLER_0_14_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ clknet_leaf_114_wb_clk_i _02317_ _00877_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08982__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16579_ clknet_leaf_124_wb_clk_i _02248_ _00808_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09120_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09379__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09051_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ _03599_ _03609_ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__and3b_2
XFILLER_0_143_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold501 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\] vssd1 vssd1
+ vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold512 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\] vssd1 vssd1
+ vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13188__X _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\] vssd1 vssd1
+ vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\] vssd1 vssd1
+ vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold545 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\] vssd1 vssd1
+ vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\] vssd1 vssd1
+ vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold567 net135 vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
X_17316__1372 vssd1 vssd1 vccd1 vccd1 _17316__1372/HI net1372 sky130_fd_sc_hd__conb_1
XFILLER_0_25_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold578 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\] vssd1 vssd1
+ vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net638 _04275_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or2_1
XANTENNA__08222__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold589 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\] vssd1 vssd1
+ vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_115_Left_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12252__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09526__B2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__mux2_1
X_09884_ _05485_ _05489_ _05494_ _04532_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout1107_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1201 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\] vssd1 vssd1
+ vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 team_04_WB.ADDR_START_VAL_REG\[10\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09842__A _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1223 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] vssd1 vssd1
+ vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
X_08835_ _03662_ _04442_ _04443_ _04444_ _04445_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a32o_1
XFILLER_0_100_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12679__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ net773 _04376_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09053__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08697_ _04304_ _04305_ _04306_ _04307_ net789 net809 vssd1 vssd1 vccd1 vccd1 _04308_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11636__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout355_X net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08892__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout522_X net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1264_X net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12597__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09318_ net777 _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09289__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1096 net1054 vssd1 vssd1 vccd1
+ vccd1 _06132_ sky130_fd_sc_hd__and3_1
XANTENNA__12061__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__mux2_1
XANTENNA__08360__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12260_ net258 net675 vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__and2_1
XANTENNA__13010__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _06271_ _06699_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_101_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_160_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12191_ _07349_ net648 vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11142_ _06216_ _06220_ net562 vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__mux2_1
XANTENNA__08132__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15950_ clknet_leaf_46_wb_clk_i _01627_ _00177_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11073_ net536 _06527_ _06561_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__and3_1
XANTENNA__08999__A1_N net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A DAT_I[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _05581_ _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and2_1
X_14901_ net1211 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__inv_2
X_15881_ clknet_leaf_73_wb_clk_i _01558_ _00108_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10898__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14832_ net1165 vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_172_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_172_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_101_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14763_ net1161 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11975_ _05736_ _05738_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16502_ clknet_leaf_11_wb_clk_i _02171_ _00731_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\]
+ sky130_fd_sc_hd__dfrtp_1
X_13714_ net993 _03101_ _03104_ net991 vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10926_ _06407_ _06413_ _06406_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__o21ai_1
X_14694_ net1104 vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ clknet_leaf_181_wb_clk_i _02102_ _00662_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\]
+ sky130_fd_sc_hd__dfrtp_1
X_13645_ _03540_ _03035_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__nand2_1
X_10857_ _06340_ _06344_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13213__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_140_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16364_ clknet_leaf_102_wb_clk_i _02033_ _00593_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13576_ _02959_ _02964_ team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1
+ _02967_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12052__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10788_ net583 _06251_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12337__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15315_ net1232 vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12527_ net2067 _07283_ net421 vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16295_ clknet_leaf_164_wb_clk_i _01964_ _00524_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13001__A1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15246_ net1204 vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__inv_2
XANTENNA__08390__X _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ net600 net237 net680 vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08103__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _06271_ _06621_ _06897_ _06277_ _06892_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__a221o_1
X_15177_ net1134 vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12389_ net222 net2584 net497 vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11563__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ team_04_WB.MEM_SIZE_REG_REG\[27\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[27\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__o221a_1
XANTENNA__12072__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14059_ net28 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1
+ vccd1 vccd1 _01527_ sky130_fd_sc_hd__o22a_1
XANTENNA__08977__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12512__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08620_ net727 _04230_ net712 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__o21a_1
XANTENNA__08278__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08482_ _04089_ _04090_ _04091_ _04092_ net784 net808 vssd1 vssd1 vccd1 vccd1 _04093_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12291__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15900__Q net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12579__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08217__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09103_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_135_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout315_A _07677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1057_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13543__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\] vssd1 vssd1
+ vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09556__B _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold331 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\] vssd1 vssd1
+ vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1224_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold342 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\] vssd1 vssd1
+ vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11554__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12751__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\] vssd1 vssd1
+ vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold364 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\] vssd1 vssd1
+ vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold375 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\] vssd1 vssd1
+ vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout800 net801 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__clkbuf_8
Xhold397 net119 vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout811 _03550_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _03721_ _03728_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and2_1
Xfanout822 _05406_ vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 net835 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__buf_4
XANTENNA__08887__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout855 net858 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__buf_4
XANTENNA__12503__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__buf_2
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout851_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _05252_ _05312_ _05475_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__or4_1
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__clkbuf_2
Xhold1020 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\] vssd1 vssd1
+ vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\] vssd1 vssd1
+ vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout899 net902 vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09380__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1042 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\] vssd1 vssd1
+ vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 net114 vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1064 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\] vssd1 vssd1
+ vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\]
+ net893 vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__mux2_1
Xhold1075 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\] vssd1 vssd1
+ vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\] vssd1 vssd1
+ vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\] vssd1 vssd1
+ vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_159_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10817__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ net701 _06190_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_159_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _03542_ _06174_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__nor2_1
XANTENNA__09511__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11490__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11691_ _06343_ _06658_ _06340_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout904_X net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12438__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13430_ _07728_ _07855_ _07730_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__a21o_1
X_10642_ net1521 team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__mux2_1
XANTENNA__08127__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12034__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13361_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] team_04_WB.MEM_SIZE_REG_REG\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[9\]
+ _06120_ net1048 vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ net1130 vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__inv_2
XANTENNA__12990__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ net2202 net499 _07600_ net438 vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a22o_1
X_13292_ _06159_ _07719_ _07721_ _07718_ net2645 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__a32o_1
XFILLER_0_122_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16080_ clknet_leaf_0_wb_clk_i _01749_ _00309_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input78_A wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ net2486 net503 _07564_ net440 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
X_15031_ net1226 vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__inv_2
XANTENNA__08097__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12173__A _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A1 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12174_ net2020 net507 _07528_ net438 vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11125_ net541 _06210_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o21ai_1
X_16982_ clknet_leaf_11_wb_clk_i _02651_ _01211_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\]
+ sky130_fd_sc_hd__dfrtp_1
X_15933_ clknet_leaf_58_wb_clk_i _01610_ _00160_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfrtp_1
X_11056_ _04440_ net544 _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__o21ai_1
X_10007_ _05606_ _05617_ _05605_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15864_ clknet_leaf_95_wb_clk_i _01541_ _00091_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_14815_ net1242 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11804__X _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14746_ net1146 vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ net691 _07129_ _07419_ net614 vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__o211a_2
XANTENNA__12273__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ net657 _06269_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__nand2_1
X_17315__1371 vssd1 vssd1 vccd1 vccd1 _17315__1371/HI net1371 sky130_fd_sc_hd__conb_1
XFILLER_0_157_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14677_ net1200 vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__inv_2
X_11889_ net687 _07360_ _07359_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16416_ clknet_leaf_137_wb_clk_i _02085_ _00645_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\]
+ sky130_fd_sc_hd__dfrtp_1
X_13628_ _07788_ _07792_ _07798_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__nor3_1
XANTENNA__13222__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11149__A1_N _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ clknet_leaf_104_wb_clk_i _02016_ _00576_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13559_ _07759_ _07821_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_763 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12981__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ clknet_leaf_14_wb_clk_i _01947_ _00507_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15229_ net1149 vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12733__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07982_ net1078 net1030 net1026 _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__or4_2
XFILLER_0_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09721_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__mux2_1
XANTENNA__08500__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _05259_ _05260_ _05261_ _05262_ net795 net803 vssd1 vssd1 vccd1 vccd1 _05263_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09901__B2 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08260__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__mux2_1
X_09583_ net580 _05192_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14738__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08534_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13461__A1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09331__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout432_A _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1174_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12016__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout220_X net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09567__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09017_ _04624_ _04625_ _04626_ _04627_ net836 net739 vssd1 vssd1 vccd1 vccd1 _04628_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout899_A net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10506__A team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1227_X net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold150 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\] vssd1 vssd1
+ vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold161 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\] vssd1 vssd1
+ vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\] vssd1 vssd1
+ vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[3\] vssd1 vssd1
+ vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\] vssd1 vssd1
+ vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13817__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _04838_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout641 _04001_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__clkbuf_2
X_09919_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\]
+ _05529_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_109_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout652 net656 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
Xfanout663 _03633_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
Xfanout674 _07554_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__buf_4
XANTENNA__08156__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout685 _07447_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__buf_4
Xfanout696 _06186_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_2
X_12930_ net241 net2573 net318 vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14324__S0 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ _07561_ net333 net389 net1930 vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14600_ net1295 vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ net704 _05827_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__o21a_1
X_15580_ net1147 vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__inv_2
XANTENNA__12255__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ net212 net2252 net322 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14531_ net1175 vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11463__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11743_ _06684_ _06861_ _07231_ _07169_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_174_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17250_ net1310 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
X_14462_ net1285 vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11674_ _03810_ net363 net360 _03809_ _07162_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ clknet_leaf_120_wb_clk_i _01870_ _00430_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\]
+ sky130_fd_sc_hd__dfrtp_1
X_13413_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__or4_1
X_17181_ clknet_leaf_90_wb_clk_i _02793_ _01410_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14393_ net1511 vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11766__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11766__B2 _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12963__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16132_ clknet_leaf_169_wb_clk_i _01801_ _00361_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11800__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] team_04_WB.MEM_SIZE_REG_REG\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__nand2_1
X_10556_ _06109_ net1563 net1020 vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07985__A3 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16063_ clknet_leaf_155_wb_clk_i _01732_ _00292_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\]
+ sky130_fd_sc_hd__dfrtp_1
X_13275_ net80 team_04_WB.ADDR_START_VAL_REG\[1\] net978 vssd1 vssd1 vccd1 vccd1 _01631_
+ sky130_fd_sc_hd__mux2_1
X_10487_ _06020_ _06055_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12715__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ net1105 vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09764__X _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ _04782_ _05279_ net822 vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__or3b_1
XFILLER_0_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12157_ _07438_ net2638 net513 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10741__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ net560 _06594_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16965_ clknet_leaf_185_wb_clk_i _02634_ _01194_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\]
+ sky130_fd_sc_hd__dfrtp_1
X_12088_ net244 net679 vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13140__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15916_ clknet_leaf_72_wb_clk_i _01593_ _00143_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11039_ net645 net550 vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nand2_1
X_16896_ clknet_leaf_137_wb_clk_i _02565_ _01125_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08242__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15847_ clknet_leaf_94_wb_clk_i _01524_ _00074_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08793__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11534__X _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15778_ net1286 vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14729_ net1133 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08250_ _03836_ _03860_ net662 vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08990__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11757__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12954__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput200 net200 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
XFILLER_0_23_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12706__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_151_Right_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12182__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10193__B1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ net778 _03575_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__nor2_1
XANTENNA__12260__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09704_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\]
+ net970 vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__mux2_1
XANTENNA__08689__A1 _04299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13682__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07896_ team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__inv_2
XANTENNA__12485__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09635_ _05242_ _05243_ _05244_ _05245_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05246_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_104_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout647_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09566_ _05173_ _05174_ _05175_ _05176_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05177_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12237__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09061__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08536__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__mux2_1
XANTENNA__13985__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09497_ _05104_ _05105_ _05106_ _05107_ net792 net812 vssd1 vssd1 vccd1 vccd1 _05108_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout814_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout435_X net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11996__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08448_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_1
XANTENNA__08861__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10089__A_N _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12945__A0 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _05611_ _05612_ _05615_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _06867_ _06868_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09728__C _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10341_ net623 _05931_ _05930_ net282 vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ net220 net2353 net304 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
X_10272_ _05536_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12011_ net247 net681 vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__and2_1
X_17314__1370 vssd1 vssd1 vccd1 vccd1 _17314__1370/HI net1370 sky130_fd_sc_hd__conb_1
XFILLER_0_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_167_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11920__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10723__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09236__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08140__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08129__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__buf_2
Xfanout471 _07668_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11067__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout482 net494 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
X_16750_ clknet_leaf_30_wb_clk_i _02419_ _00979_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13962_ net153 net1064 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__and2_1
Xfanout493 net494 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_4
X_15701_ net1258 vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_79_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12913_ _07615_ net347 net387 net2017 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a22o_1
X_16681_ clknet_leaf_122_wb_clk_i _02350_ _00910_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\]
+ sky130_fd_sc_hd__dfrtp_1
X_13893_ _03159_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15632_ net1163 vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__inv_2
X_12844_ _07542_ net337 net393 net2006 vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15563_ net1159 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12775_ _07502_ net348 net399 net2634 vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__a22o_1
X_17302_ net1358 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
X_14514_ net1192 vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__inv_2
X_11726_ _06520_ _06521_ _07199_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__nor4_1
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08663__X _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15494_ net1104 vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11451__A3 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13189__B1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ net135 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ net1277 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__inv_2
X_11657_ _04610_ _04642_ net358 _07145_ net462 vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o311a_1
XFILLER_0_153_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12936__B1 _07676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ net61 _06145_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17164_ clknet_leaf_84_wb_clk_i _02776_ _01393_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14376_ net1549 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17197__Q team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _07061_ _07076_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__xor2_1
XANTENNA__12345__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ clknet_leaf_182_wb_clk_i _01784_ _00344_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_13327_ net1086 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 _07753_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold908 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\] vssd1 vssd1
+ vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1097 net1053 vssd1 vssd1 vccd1
+ vccd1 _06098_ sky130_fd_sc_hd__and3_1
X_17095_ clknet_leaf_91_wb_clk_i _02730_ _01324_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold919 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\] vssd1 vssd1
+ vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09935__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16046_ clknet_leaf_32_wb_clk_i _01715_ _00275_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_13258_ net78 team_04_WB.ADDR_START_VAL_REG\[18\] net975 vssd1 vssd1 vccd1 vccd1
+ _01648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12164__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12209_ _07402_ net649 vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__and2_1
XANTENNA__13900__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ net1031 net1027 net1077 vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__a21oi_2
XANTENNA__10175__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15672__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16948_ clknet_leaf_1_wb_clk_i _02617_ _01177_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12467__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16879_ clknet_leaf_188_wb_clk_i _02548_ _01108_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\]
+ sky130_fd_sc_hd__dfrtp_1
X_09420_ net589 _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\]
+ net893 vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__mux2_1
XANTENNA__13967__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11978__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08302_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__mux2_1
X_09282_ _03724_ _03835_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10650__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout228_A _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08164_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14129__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08095_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12823__X _07672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload70 clknet_leaf_51_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload70/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload81 clknet_leaf_52_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__clkinv_2
Xclkload92 clknet_leaf_146_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload92/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09056__S net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _04604_ _04605_ _04606_ _04607_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04608_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout764_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__nor2_1
XANTENNA__08895__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout931_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] vssd1 vssd1
+ vccd1 vccd1 _03494_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09618_ _05225_ _05226_ _05227_ _05228_ net834 net746 vssd1 vssd1 vccd1 vccd1 _05229_
+ sky130_fd_sc_hd__mux4_1
X_10890_ _06368_ _06372_ _06378_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nor3_1
XANTENNA__11418__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__S0 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\]
+ net951 vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__mux2_1
XANTENNA__11969__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11513__S0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12091__B1 _07500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12560_ _07527_ net483 net417 net2097 vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XANTENNA__12630__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _04977_ _06248_ _06824_ _06948_ _06999_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12491_ _07488_ net488 net426 net1686 vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a22o_1
XANTENNA__12446__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11988__C _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12918__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ _03422_ net819 _03421_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__and3b_1
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_126_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11442_ net286 _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__or2_1
XANTENNA__08135__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14161_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__nor2_1
X_11373_ team_04_WB.MEM_SIZE_REG_REG\[14\] _06507_ team_04_WB.MEM_SIZE_REG_REG\[15\]
+ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_169_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07974__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input60_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10324_ _05753_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__xor2_1
X_13112_ _07544_ net371 net298 net1913 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a22o_1
X_14092_ net1448 _06130_ net1035 vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10255_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] net1055 _05853_
+ _05855_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13043_ _07504_ net375 net306 net1971 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__a22o_1
XANTENNA__12181__A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12697__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1200 net1201 vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_4
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] net1055 _05792_
+ _05794_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
Xfanout1222 net1224 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__buf_2
Xfanout1233 net1234 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
Xfanout1244 net1252 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__buf_4
Xfanout1255 net1257 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__buf_4
X_16802_ clknet_leaf_146_wb_clk_i _02471_ _01031_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1266 net1280 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__buf_2
Xfanout1277 net1278 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__buf_4
X_14994_ net1236 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__inv_2
XANTENNA__12449__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1288 net1297 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__buf_2
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
X_16733_ clknet_leaf_131_wb_clk_i _02402_ _00962_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\]
+ sky130_fd_sc_hd__dfrtp_1
X_13945_ team_04_WB.ADDR_START_VAL_REG\[0\] _03078_ net1040 vssd1 vssd1 vccd1 vccd1
+ _03305_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13216__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload6_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16664_ clknet_leaf_149_wb_clk_i _02333_ _00893_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\]
+ sky130_fd_sc_hd__dfrtp_1
X_13876_ _02941_ _03258_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ net1270 vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12827_ _07525_ net341 net392 net1855 vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16595_ clknet_leaf_183_wb_clk_i _02264_ _00824_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ net1151 vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08393__X _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ _07485_ net334 net397 net2122 vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12621__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11709_ _07185_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15477_ net1209 vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12689_ _06189_ _07665_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__or2_4
XANTENNA__11260__A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17216_ net1422 _02826_ _01459_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12909__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ net1289 vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__inv_2
XANTENNA__09001__Y _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_96_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17147_ clknet_leaf_85_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[1\]
+ _01376_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14359_ net1262 vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold705 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\] vssd1 vssd1
+ vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold716 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\] vssd1 vssd1
+ vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold727 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\] vssd1 vssd1
+ vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14126__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold738 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\] vssd1 vssd1
+ vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17078_ clknet_leaf_45_wb_clk_i _00026_ _01307_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold749 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\] vssd1 vssd1
+ vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08920_ _04359_ _04414_ _04477_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16029_ clknet_leaf_129_wb_clk_i _01698_ _00258_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10604__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13885__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08851_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13637__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\]
+ net866 vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__mux2_1
XANTENNA__09604__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__B net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12860__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09403_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14062__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ _04941_ _04942_ _04943_ _04944_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04945_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12612__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09265_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\]
+ net925 vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout512_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12266__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1254_A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _03823_ _03824_ _03825_ _03826_ net791 net812 vssd1 vssd1 vccd1 vccd1 _03827_
+ sky130_fd_sc_hd__mux4_1
X_09196_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08044__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14117__A2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload170 clknet_leaf_83_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload170/Y sky130_fd_sc_hd__inv_6
X_08078_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout881_A net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout979_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10040_ _05555_ _05650_ _05554_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09862__X _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__C net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11329__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\] vssd1 vssd1
+ vccd1 vccd1 net1447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 net169 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold76 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\] vssd1 vssd1 vccd1
+ vccd1 net1513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[24\] vssd1 vssd1
+ vccd1 vccd1 net1524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[8\]
+ vssd1 vssd1 vccd1 vccd1 net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _04782_ _05280_ net822 vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__or3b_2
XANTENNA__12300__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13730_ _03118_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10942_ net632 _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12851__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ net995 _03047_ _03051_ _07691_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__a22o_1
X_10873_ _04556_ _06360_ _06361_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__and3_1
XANTENNA__14053__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14656__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ net1116 vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__inv_2
X_12612_ _07581_ net488 net414 net1958 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11999__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16380_ clknet_leaf_128_wb_clk_i _02049_ _00609_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09155__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ _06973_ net271 net710 vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_130_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12603__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ net1168 vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__inv_2
X_12543_ net2123 net253 net420 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08902__S1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08283__A2 _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15262_ net1215 vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12474_ net608 net233 net683 vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17001_ clknet_leaf_100_wb_clk_i _02670_ _01230_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\]
+ sky130_fd_sc_hd__dfrtp_1
X_14213_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ _03412_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__or2_1
X_11425_ _06633_ _06913_ net581 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__a21oi_1
X_15193_ net1246 vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__inv_2
XANTENNA_7 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14108__A2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14144_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03356_
+ _03362_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__or3_1
X_11356_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__inv_2
XANTENNA__12119__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _05578_ _05580_ _05635_ net623 _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__o311a_1
X_14075_ net1492 _06096_ net1035 vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__mux2_1
X_11287_ net576 _06702_ _06769_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_94_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13026_ _07487_ net376 net308 net1654 vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__a22o_1
X_10238_ _05563_ _05644_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1030 _03538_ vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13735__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10169_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] net1056 _05545_
+ _05779_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a22o_1
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_2
Xfanout1063 _03350_ vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13619__B2 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1074 net1076 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09424__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1085 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 net1085 sky130_fd_sc_hd__buf_2
Xfanout1096 net1097 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_2
X_14977_ net1150 vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__inv_2
XANTENNA__13095__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ net1827 net1071 net1040 _03295_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__a22o_1
X_16716_ clknet_leaf_112_wb_clk_i _02385_ _00945_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12842__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16647_ clknet_leaf_24_wb_clk_i _02316_ _00876_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\]
+ sky130_fd_sc_hd__dfrtp_1
X_13859_ _02873_ _03226_ _03229_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_174_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14044__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16578_ clknet_leaf_147_wb_clk_i _02247_ _00807_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__Y _06750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15529_ net1134 vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12086__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ _04657_ _04658_ _04659_ _04660_ net786 net806 vssd1 vssd1 vccd1 vccd1 _04661_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08001_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__or2_2
XFILLER_0_128_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold502 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\] vssd1 vssd1
+ vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\] vssd1 vssd1
+ vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\] vssd1 vssd1
+ vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold535 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\] vssd1 vssd1
+ vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold546 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\] vssd1 vssd1
+ vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\] vssd1 vssd1
+ vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\] vssd1 vssd1
+ vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ net592 _04167_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__xnor2_1
Xhold579 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\] vssd1 vssd1
+ vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08903_ net728 _04513_ net712 vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__o21a_1
X_09883_ _05491_ _05493_ _04755_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_148_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09082__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1202 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\] vssd1 vssd1
+ vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\] _03650_ _03652_
+ _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o311a_1
Xhold1213 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] vssd1 vssd1
+ vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1224 team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1002_A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _04372_ _04373_ _04374_ _04375_ net789 net810 vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_174_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout462_A _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11097__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08696_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__mux2_1
XANTENNA__12833__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14476__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14035__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09317_ _04924_ _04925_ _04926_ _04927_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04928_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_118_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10509__A team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08896__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1257_X net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09248_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09509__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ net562 _06240_ _06612_ _06698_ _06246_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__a32o_1
X_12190_ net2034 net509 _07536_ net459 vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a22o_1
XANTENNA__09765__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ _06328_ _06629_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11072_ net664 _05374_ _05343_ _03834_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__a211o_2
XFILLER_0_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput100 wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11324__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _05585_ _05631_ _05586_ _05584_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o211ai_1
X_14900_ net1214 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__inv_2
X_15880_ clknet_leaf_79_wb_clk_i _01557_ _00107_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08820__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09244__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A DAT_I[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14831_ net1199 vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14762_ net1124 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__inv_2
XANTENNA__08489__C1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11974_ net2210 net528 net455 _07433_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a22o_1
XANTENNA__12824__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ clknet_leaf_35_wb_clk_i _02170_ _00730_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13713_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _05934_ net1102
+ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10925_ _06407_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14693_ net1113 vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16432_ clknet_leaf_1_wb_clk_i _02101_ _00661_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\]
+ sky130_fd_sc_hd__dfrtp_1
X_13644_ net993 _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_141_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10856_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16363_ clknet_leaf_25_wb_clk_i _02032_ _00592_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\]
+ sky130_fd_sc_hd__dfrtp_1
X_13575_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ net645 _06269_ _06270_ _06275_ _06260_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__o311a_1
X_15314_ net1244 vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__inv_2
X_12526_ net2251 net218 net420 vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__mux2_1
X_16294_ clknet_leaf_17_wb_clk_i _01963_ _00523_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15245_ net1199 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ net2444 net428 _07648_ net520 vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10706__X _06195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15010__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11408_ _06845_ _06896_ net576 vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__mux2_1
XANTENNA__09419__S net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09300__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15176_ net1125 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__inv_2
X_12388_ net229 net2513 net497 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__mux2_1
XANTENNA__12353__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11563__A2 _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ team_04_WB.MEM_SIZE_REG_REG\[26\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[26\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_91_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11339_ net553 _06827_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09943__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ net29 net1063 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1
+ vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
X_13009_ net606 _07469_ net471 net311 net1790 vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15680__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
XANTENNA__08993__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08581__X _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13199__X _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ _04610_ _04642_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold310 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\] vssd1 vssd1
+ vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08233__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold321 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\] vssd1 vssd1
+ vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\] vssd1 vssd1
+ vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\] vssd1 vssd1
+ vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\] vssd1 vssd1
+ vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_159_72 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold365 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\] vssd1 vssd1
+ vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\] vssd1 vssd1
+ vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold387 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\] vssd1 vssd1
+ vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout801 net804 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_8
Xhold398 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\] vssd1 vssd1
+ vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ _03721_ _03728_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nor2_1
Xfanout812 net815 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
Xfanout823 net830 vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_4
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__buf_4
XANTENNA__09055__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12503__A1 _07500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_A _07482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net858 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__clkbuf_4
X_09866_ _05378_ net533 _05404_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__a21boi_1
Xfanout867 net871 vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 net883 vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__buf_4
Xhold1010 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\] vssd1 vssd1
+ vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\] vssd1 vssd1
+ vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 net895 vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09064__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
Xhold1032 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\] vssd1 vssd1
+ vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\] vssd1 vssd1
+ vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _05405_ _05407_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__or2_1
Xhold1054 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\] vssd1 vssd1
+ vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\] vssd1 vssd1
+ vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1076 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\] vssd1 vssd1
+ vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08748_ _04328_ _04357_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__xnor2_1
Xhold1087 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\] vssd1 vssd1
+ vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\] vssd1 vssd1
+ vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_2_0_wb_clk_i_X clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10710_ _04726_ _05444_ _03635_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__o21a_1
X_11690_ net286 _07175_ _07176_ _07178_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__or4_2
XFILLER_0_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ net1508 team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_923 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13360_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\] team_04_WB.MEM_SIZE_REG_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10572_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06120_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_165_Right_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12990__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ net239 net668 vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13291_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\] _07720_
+ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12454__A net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15030_ net1223 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__inv_2
XANTENNA__09239__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ net241 net672 vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09294__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12173__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ _07289_ net647 vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__and2_1
XANTENNA__10753__A0 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ net532 _06214_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16981_ clknet_leaf_12_wb_clk_i _02650_ _01210_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\]
+ sky130_fd_sc_hd__dfrtp_1
X_15932_ clknet_leaf_58_wb_clk_i _01609_ _00159_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfrtp_1
X_11055_ net591 net544 vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10006_ _05609_ _05616_ _05608_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__a21oi_1
X_15863_ clknet_leaf_94_wb_clk_i _01540_ _00090_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10421__B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14814_ net1217 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09702__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745_ net1235 vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__inv_2
X_11957_ _07398_ _07418_ _07417_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_28_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13224__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11533__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15005__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ net580 _06394_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__nor2_1
XANTENNA__11481__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14676_ net1225 vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__inv_2
X_11888_ team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07360_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16415_ clknet_leaf_161_wb_clk_i _02084_ _00644_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\]
+ sky130_fd_sc_hd__dfrtp_1
X_13627_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10839_ _03892_ _06325_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16346_ clknet_leaf_39_wb_clk_i _02015_ _00575_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09938__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ _06880_ net273 vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12981__A1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12509_ _07506_ net480 net424 net1803 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ clknet_leaf_33_wb_clk_i _01946_ _00506_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\]
+ sky130_fd_sc_hd__dfrtp_1
X_13489_ net996 _02879_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15228_ net1130 vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15159_ net1230 vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__inv_2
XANTENNA__08988__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07981_ team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] team_04_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09720_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\]
+ net968 vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__mux2_1
XANTENNA__11708__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12497__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08289__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__mux2_1
XANTENNA__09901__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08260__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08533_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__mux2_1
XANTENNA__13997__B1 _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11443__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08464_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\]
+ net853 vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__mux2_1
XANTENNA__08228__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12258__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08395_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14754__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_A _07656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1167_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12421__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07979__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09200__X _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12972__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12274__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09016_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout794_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13921__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold151 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold162 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[5\] vssd1 vssd1
+ vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08898__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\] vssd1 vssd1
+ vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09583__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\] vssd1 vssd1
+ vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\] vssd1 vssd1
+ vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09028__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net621 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
Xfanout631 _04838_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_2
X_09918_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _05528_ vssd1
+ vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout653 net655 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XANTENNA__12488__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08199__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08156__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout664 net665 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 _07554_ vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
Xfanout686 net688 vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
Xfanout697 _06184_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__clkbuf_4
X_09849_ _05458_ _05459_ _05451_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__o21ba_2
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12860_ _07560_ net341 net388 net2158 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__a22o_1
XANTENNA__14324__S1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11811_ net686 _07292_ _07291_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__a21oi_1
X_12791_ net211 net2415 net323 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ net1173 vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11742_ _06732_ _06818_ _06881_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__or4_1
XFILLER_0_138_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12660__A0 _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08138__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ net1186 vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ net644 _03808_ net359 vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16200_ clknet_leaf_112_wb_clk_i _01869_ _00429_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\]
+ sky130_fd_sc_hd__dfrtp_1
X_13412_ team_04_WB.MEM_SIZE_REG_REG\[20\] _07831_ _07837_ vssd1 vssd1 vccd1 vccd1
+ _07838_ sky130_fd_sc_hd__a21o_1
XANTENNA__07977__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input90_A wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__or4b_1
X_17180_ clknet_leaf_91_wb_clk_i _02792_ _01409_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12412__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14392_ net1513 vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_133_Left_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12963__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16131_ clknet_leaf_117_wb_clk_i _01800_ _00360_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_13343_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] team_04_WB.MEM_SIZE_REG_REG\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__xor2_2
XFILLER_0_148_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11800__B net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10555_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[15\]
+ _06108_ net1047 vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16062_ clknet_leaf_143_wb_clk_i _01731_ _00291_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_13274_ net91 team_04_WB.ADDR_START_VAL_REG\[2\] net978 vssd1 vssd1 vccd1 vccd1 _01632_
+ sky130_fd_sc_hd__mux2_1
X_10486_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] net1006 _06061_ _06062_
+ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15013_ net1109 vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _04783_ _05280_ net822 vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__and3_4
XANTENNA__10726__A0 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11923__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ net222 net2622 net513 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__mux2_1
XANTENNA__08601__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10703__Y _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13219__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ net531 _06262_ _06595_ net557 vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__o211a_1
X_12087_ net2180 net353 _07498_ net447 vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16964_ clknet_leaf_167_wb_clk_i _02633_ _01193_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_142_Left_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15915_ clknet_leaf_72_wb_clk_i _01592_ _00142_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ _03721_ net544 vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nand2_1
XANTENNA__11151__A0 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08242__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16895_ clknet_leaf_157_wb_clk_i _02564_ _01124_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ clknet_leaf_98_wb_clk_i _01523_ _00073_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_15777_ net1286 vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__inv_2
X_12989_ net699 _07448_ _07666_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_82_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14728_ net1117 vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__inv_2
XANTENNA__12651__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12078__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ net1182 vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__inv_2
XANTENNA__12793__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14574__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11550__X _07039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12403__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11757__A2 _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11710__B _06592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16329_ clknet_leaf_102_wb_clk_i _01998_ _00558_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput201 net201 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_0_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12182__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10193__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_160_Left_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07964_ _03571_ _03572_ _03573_ _03574_ net787 net810 vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_147_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09703_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\]
+ net966 vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__mux2_1
XANTENNA__10061__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09886__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07895_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1 _03510_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout375_A _07679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__mux2_1
XANTENNA__14101__X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08747__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09565_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout542_A _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1284_A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08516_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12642__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__mux2_1
XANTENNA__11996__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout330_X net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11901__A net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ net770 _03982_ net761 vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09497__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10340_ _05627_ _05929_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10271_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _05535_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\]
+ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09517__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ net2515 net515 _07458_ net438 vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_143_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08421__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08129__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout450 net452 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_4
Xfanout461 _07252_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_2
Xfanout472 net473 vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
X_13961_ _03973_ net262 net598 _03314_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a31o_1
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout494 _07655_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_6
XANTENNA__13673__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__B2 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15700_ net1262 vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__inv_2
X_12912_ _07614_ net330 net384 net1905 vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22o_1
X_16680_ clknet_leaf_114_wb_clk_i _02349_ _00909_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\]
+ sky130_fd_sc_hd__dfrtp_1
X_13892_ _03168_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__or2_1
XANTENNA__12881__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09252__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15631_ net1195 vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__inv_2
X_12843_ _07541_ net338 net393 net2021 vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11083__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15562_ net1105 vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12774_ _07501_ net350 net399 net1850 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a22o_1
XANTENNA__12633__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17301_ net1357 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
X_14513_ net1191 vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11725_ _06628_ _07184_ _07200_ _07213_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__or4b_1
XFILLER_0_138_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15493_ net1109 vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__inv_2
XANTENNA__11159__A_N _06227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17232_ net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input93_X net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ net1277 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11656_ _04610_ _04642_ net361 vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ _06142_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__nor2_2
X_17163_ clknet_leaf_84_wb_clk_i _02775_ _01392_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_86_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14375_ net1561 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11587_ net708 _07075_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ clknet_leaf_7_wb_clk_i _01783_ _00343_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_13326_ net1085 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 _07752_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_101_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10538_ _06097_ net1577 net1022 vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__mux2_1
X_17094_ clknet_leaf_91_wb_clk_i _02729_ _01323_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold909 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\] vssd1 vssd1
+ vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16045_ clknet_leaf_43_wb_clk_i _01714_ _00274_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_13257_ net79 team_04_WB.ADDR_START_VAL_REG\[19\] net975 vssd1 vssd1 vccd1 vccd1
+ _01649_ sky130_fd_sc_hd__mux2_1
XANTENNA__13738__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _06006_ _06013_ _06047_ _03528_ _03513_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__o32ai_1
XANTENNA__09935__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09427__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12164__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12208_ net2336 net510 _07545_ net458 vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13188_ net1031 net1027 net1077 vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__a21o_2
XANTENNA__10175__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11911__A2 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _07327_ net2582 net512 vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09951__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16947_ clknet_leaf_181_wb_clk_i _02616_ _01176_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14569__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16878_ clknet_leaf_27_wb_clk_i _02547_ _01107_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12872__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15829_ clknet_leaf_93_wb_clk_i _01506_ _00056_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\]
+ net893 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__mux2_1
XANTENNA__12624__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13967__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08301_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ net766 _04891_ _04880_ _04874_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08232_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__mux2_1
XANTENNA__10650__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08163_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\]
+ net946 vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux2_1
XANTENNA__14129__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\]
+ net919 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10056__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload60 clknet_leaf_37_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_6
Xclkload71 clknet_leaf_53_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_77_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload82 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__inv_4
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1032_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload93 clknet_leaf_147_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload93/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_149_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08241__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout492_A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09861__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _03556_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13655__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09859__B2 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07878_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 _03493_ sky130_fd_sc_hd__inv_2
XANTENNA__12863__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14198__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout924_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ _05155_ _05156_ _05157_ _05158_ net795 net813 vssd1 vssd1 vccd1 vccd1 _05159_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12615__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_120_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09800__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09479_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12091__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11510_ _04976_ _06253_ _06257_ _04975_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_163_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12490_ _07487_ net487 net426 net1738 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__a22o_1
XANTENNA__08416__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12918__A1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11441_ _06924_ _06927_ _06929_ _06925_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__or4b_1
XFILLER_0_110_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13040__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14160_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nor2_1
XANTENNA__11051__C1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ _06858_ _06860_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13111_ _07543_ net367 net298 net1705 vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_169_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10323_ _05704_ _05705_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14091_ net1459 _06128_ net1034 vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__mux2_1
XANTENNA__14135__A3 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_166_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_166_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09247__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input53_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _07503_ net380 net309 net1787 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__a22o_1
X_10254_ net277 _05854_ net1074 vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__o21a_1
XANTENNA__08151__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12181__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__clkbuf_4
Xfanout1212 net1220 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__buf_4
X_10185_ net278 _05793_ net1074 vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__o21a_1
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__buf_4
XFILLER_0_100_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1234 net1253 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__clkbuf_2
X_16801_ clknet_leaf_133_wb_clk_i _02470_ _01030_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1245 net1252 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__buf_2
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_2
Xfanout1267 net1269 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13646__A2 _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _05523_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_4
Xfanout1278 net1279 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__buf_2
X_14993_ net1266 vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__inv_2
Xfanout291 _07684_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_4
Xfanout1289 net1293 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__buf_4
XANTENNA__11657__A1 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ clknet_leaf_127_wb_clk_i _02401_ _00961_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\]
+ sky130_fd_sc_hd__dfrtp_1
X_13944_ _03081_ net1040 _03304_ net1071 net2490 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a32o_1
XANTENNA__12854__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13875_ _03194_ _03198_ _02943_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__a21oi_1
X_16663_ clknet_leaf_174_wb_clk_i _02332_ _00892_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12826_ _07524_ net341 net394 net1615 vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__a22o_1
X_15614_ net1216 vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__inv_2
XANTENNA__12606__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16594_ clknet_leaf_7_wb_clk_i _02263_ _00823_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09710__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15545_ net1248 vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__inv_2
X_12757_ net701 _07483_ _07663_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__or3_4
XFILLER_0_16_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13232__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ net706 _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15476_ net1235 vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ net614 _06196_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12909__A1 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17215_ net1421 _02825_ _01457_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_14427_ net1289 vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13031__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11639_ _06206_ _07121_ _07127_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__nor3_1
XANTENNA__14852__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17146_ clknet_leaf_85_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[0\]
+ _01375_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14358_ net1262 vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09946__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\] vssd1 vssd1
+ vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold717 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\] vssd1 vssd1
+ vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11593__B1 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13309_ net1083 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 _07735_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_141_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold728 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\] vssd1 vssd1
+ vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10591__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17077_ clknet_leaf_45_wb_clk_i _00025_ _01306_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14289_ _03458_ _03459_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__nor2_1
Xhold739 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\] vssd1 vssd1
+ vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16028_ clknet_leaf_129_wb_clk_i _01697_ _00257_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10604__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08850_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__mux2_1
XANTENNA__11896__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08996__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _04388_ _04389_ _04390_ _04391_ net827 net743 vssd1 vssd1 vccd1 vccd1 _04392_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13098__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12845__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09402_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13619__A2_N net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09333_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__mux2_1
XANTENNA__13270__A0 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_wb_clk_i_X clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12073__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_A _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09264_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\]
+ net925 vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12266__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__mux2_1
XANTENNA__13022__B1 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout505_A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1247_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09856__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\]
+ net924 vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08044__A3 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08077_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12282__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload160 clknet_leaf_103_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload160/Y sky130_fd_sc_hd__inv_6
Xclkload171 clknet_leaf_84_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload171/Y sky130_fd_sc_hd__bufinv_16
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_692 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13325__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11887__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1202_X net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\] vssd1 vssd1 vccd1
+ vccd1 net1470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08979_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__mux2_1
Xhold55 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[21\]
+ vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10530__A team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold88 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[23\] vssd1 vssd1
+ vccd1 vccd1 net1525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12836__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14002__A _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11990_ _04783_ _05279_ net822 vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__and3_1
Xhold99 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[17\]
+ vssd1 vssd1 vccd1 vccd1 net1536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12300__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _04812_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _03026_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__or2_1
X_10872_ _06358_ _06359_ _04585_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12611_ _07580_ net492 net414 net2367 vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13591_ _02980_ _02981_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15330_ net1219 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__inv_2
X_12542_ net2047 net254 net421 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__mux2_1
XANTENNA__11811__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15261_ net1147 vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__inv_2
XANTENNA__11080__B _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ net523 net607 _07474_ net430 net1750 vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a32o_1
XANTENNA__13013__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14212_ _03365_ _03413_ _03414_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[5\]
+ sky130_fd_sc_hd__and3_1
X_17000_ clknet_leaf_114_wb_clk_i _02669_ _01229_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13564__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ net574 _06911_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15192_ net1206 vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__inv_2
XANTENNA__08670__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] _03363_
+ team_04_WB.instance_to_wrap.final_design.h_out vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _06689_ _06765_ net558 vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12119__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _05578_ _05580_ _05635_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__o21ai_1
X_14074_ net1478 _06094_ net1032 vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11286_ net289 _06771_ _06773_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a22o_1
X_13025_ _07486_ net371 net308 net1612 vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22o_1
X_10237_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] net1074 _05839_
+ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__o21ba_1
Xfanout1020 _06073_ vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__clkbuf_4
Xfanout1031 _03538_ vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09705__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1042 _03244_ vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__clkbuf_4
Xfanout1053 net1054 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
X_10168_ net622 _05661_ _05778_ net281 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a211o_1
Xfanout1064 net1065 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__buf_2
XANTENNA__13227__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1075 net1076 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_2
Xfanout1086 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\] vssd1 vssd1 vccd1
+ vccd1 net1086 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15008__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12827__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12131__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _04786_ vssd1
+ vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__nand2_1
X_14976_ net1220 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_63_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16715_ clknet_leaf_31_wb_clk_i _02384_ _00944_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\]
+ sky130_fd_sc_hd__dfrtp_1
X_13927_ _03098_ _03141_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16646_ clknet_leaf_17_wb_clk_i _02315_ _00875_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\]
+ sky130_fd_sc_hd__dfrtp_1
X_13858_ _02873_ _03226_ _03229_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__or3_1
XFILLER_0_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09440__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ net255 net2272 net325 vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16577_ clknet_leaf_134_wb_clk_i _02246_ _00806_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\]
+ sky130_fd_sc_hd__dfrtp_1
X_13789_ _03171_ _03175_ _03178_ team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1
+ vccd1 _03180_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_174_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ net1116 vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12086__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13004__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ net1172 vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08000_ net1078 net1031 net1027 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_96_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12358__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\] vssd1 vssd1
+ vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17129_ clknet_leaf_75_wb_clk_i net1499 _01358_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold514 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\] vssd1 vssd1
+ vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold525 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\] vssd1 vssd1
+ vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold547 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\] vssd1 vssd1
+ vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ net594 _04114_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__and2_1
Xhold558 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\] vssd1 vssd1
+ vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\] vssd1 vssd1
+ vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09606__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08902_ _04509_ _04510_ _04511_ _04512_ net829 net736 vssd1 vssd1 vccd1 vccd1 _04513_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09882_ _04868_ _05490_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09082__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08833_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__or3_1
Xhold1203 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\] vssd1 vssd1
+ vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] vssd1
+ vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09842__C _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1225 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12818__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11097__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout455_A net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08593__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1197_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Right_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09350__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12046__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_X net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09316_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__mux2_1
XANTENNA__12597__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13794__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08896__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout410_X net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13546__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_147 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13010__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ net728 _03739_ net714 vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08973__A1 _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _06331_ _06487_ _06330_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13836__A team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _06557_ _06559_ net536 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__mux2_1
Xinput101 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_1
X_10022_ _05583_ _05632_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__nor2_1
XANTENNA__09525__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ net1200 vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__inv_2
XANTENNA__12809__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input16_A DAT_I[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ net1136 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__inv_2
X_11973_ net654 net221 vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12285__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ clknet_leaf_2_wb_clk_i _02169_ _00729_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\]
+ sky130_fd_sc_hd__dfrtp_1
X_13712_ net999 _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__or2_1
X_10924_ _05379_ _06411_ _06410_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__a21oi_1
X_14692_ net1171 vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14026__A2 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13234__A0 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16431_ clknet_leaf_187_wb_clk_i _02100_ _00660_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\]
+ sky130_fd_sc_hd__dfrtp_1
X_13643_ _07798_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__or2_1
X_10855_ _04166_ _06341_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12187__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12588__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13574_ team_04_WB.ADDR_START_VAL_REG\[14\] _02959_ _02964_ vssd1 vssd1 vccd1 vccd1
+ _02965_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16362_ clknet_leaf_163_wb_clk_i _02031_ _00591_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10786_ net567 _06239_ _06271_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ net2183 net220 net422 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__mux2_1
X_15313_ net1270 vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16293_ clknet_leaf_20_wb_clk_i _01962_ _00522_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_181_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_181_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_48_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13537__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ net602 net248 net680 vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15244_ net1121 vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__inv_2
XANTENNA__08604__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13001__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ net555 _06767_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__a21oi_1
X_15175_ net1139 vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12387_ net231 net2338 net497 vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__mux2_1
X_14126_ team_04_WB.MEM_SIZE_REG_REG\[25\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[25\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__o221a_1
XANTENNA__10220__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12760__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ _06552_ _06557_ net536 vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11563__A3 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14057_ net30 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1
+ vccd1 vccd1 _01529_ sky130_fd_sc_hd__o22a_1
X_11269_ net706 _06734_ net284 vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__or3_2
XANTENNA__09943__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12512__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ net610 _07468_ net473 net312 net1778 vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a32o_1
XFILLER_0_158_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14959_ net1141 vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__inv_2
XANTENNA__12796__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14017__A2 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13225__A0 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16629_ clknet_leaf_33_wb_clk_i _02298_ _00858_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12028__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12579__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09032_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__inv_2
XANTENNA__15201__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11539__A0 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold300 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\] vssd1 vssd1
+ vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\] vssd1 vssd1
+ vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12200__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\] vssd1 vssd1
+ vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\] vssd1 vssd1
+ vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12751__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\] vssd1 vssd1
+ vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\] vssd1 vssd1
+ vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold366 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\] vssd1 vssd1
+ vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10064__B _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold377 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\] vssd1 vssd1
+ vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\] vssd1 vssd1
+ vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net803 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__clkbuf_8
X_09934_ net277 _05544_ net1074 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__o21a_1
Xhold399 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\] vssd1 vssd1
+ vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09853__B net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout813 net815 vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__buf_4
Xfanout824 net830 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
XANTENNA__09055__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout835 net838 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09345__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout846 net859 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12503__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input8_A DAT_I[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout857 net858 vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_4
X_09865_ _05378_ net532 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__and2_1
Xhold1000 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\] vssd1 vssd1
+ vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net870 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__clkbuf_4
Xhold1011 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\] vssd1 vssd1
+ vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net880 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09380__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1022 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\] vssd1 vssd1
+ vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\] vssd1 vssd1
+ vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
X_09796_ _03637_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__and2_1
Xhold1044 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\] vssd1 vssd1
+ vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1055 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\] vssd1 vssd1
+ vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\] vssd1 vssd1
+ vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _04328_ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__and2_1
Xhold1077 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\] vssd1 vssd1
+ vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\] vssd1 vssd1
+ vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1099 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\] vssd1 vssd1
+ vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout837_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10278__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08678_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_159_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ net1498 team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _06119_ net1539 net1021 vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XANTENNA__12294__X _07591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ net2328 net499 _07599_ net440 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\] vssd1 vssd1 vccd1
+ vccd1 _07720_ sky130_fd_sc_hd__and3_1
XANTENNA__08424__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ net2290 net503 _07563_ net438 vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__a22o_1
XANTENNA__09294__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12742__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ net2081 net508 _07527_ net445 vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__a22o_1
XANTENNA__10753__A1 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13566__A team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11123_ net533 _06212_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_1
X_16980_ clknet_leaf_1_wb_clk_i _02649_ _01209_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ clknet_leaf_58_wb_clk_i _01608_ _00158_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfrtp_1
X_11054_ net636 _04557_ net550 vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__mux2_1
XANTENNA__11702__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _05612_ _05615_ _05611_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__a21o_1
X_15862_ clknet_leaf_94_wb_clk_i _01539_ _00089_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_14813_ net1149 vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11814__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ net1208 vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__inv_2
X_11956_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[4\] team_04_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ net266 vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ net580 _06394_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11887_ net705 _05907_ _07358_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__o21ai_1
X_14675_ net1227 vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__inv_2
XANTENNA__13758__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ clknet_leaf_158_wb_clk_i _02083_ _00643_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13626_ _03015_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10838_ _03891_ _06325_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11769__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11820__Y _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16345_ clknet_leaf_177_wb_clk_i _02014_ _00574_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\]
+ sky130_fd_sc_hd__dfrtp_1
X_13557_ _02944_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__nor2_1
XANTENNA__09938__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _05450_ _05464_ _05470_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13240__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07988__A2 _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12981__A2 _07403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ _07505_ net485 net425 net1810 vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a22o_1
X_13488_ net1092 _02878_ net1043 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__o2bb2a_1
X_16276_ clknet_leaf_4_wb_clk_i _01945_ _00505_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10992__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15227_ net1113 vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__inv_2
X_12439_ net2233 net435 _07640_ net525 vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09954__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ net1221 vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11548__X _07037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ team_04_WB.MEM_SIZE_REG_REG\[8\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[8\]
+ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__a22o_2
XFILLER_0_10_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14071__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1009 _03590_ vssd1 vssd1 vccd1
+ vccd1 _03591_ sky130_fd_sc_hd__a21o_1
X_15089_ net1266 vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09165__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09362__A1 _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__mux2_1
X_09581_ _05167_ _05191_ net664 vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__mux2_2
XANTENNA__12249__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13513__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08548__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08463_ _04070_ _04071_ _04072_ _04073_ net825 net734 vssd1 vssd1 vccd1 vccd1 _04074_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10059__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_154_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12421__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout320_A net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08244__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_171_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12274__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__mux2_1
XANTENNA__10506__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07936__X _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\] vssd1 vssd1
+ vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[12\] vssd1
+ vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold152 team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] vssd1
+ vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout787_A net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\] vssd1 vssd1
+ vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold174 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\] vssd1 vssd1
+ vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\] vssd1 vssd1
+ vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10803__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\] vssd1 vssd1
+ vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09028__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout610 net612 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
Xfanout621 net624 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09075__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\]
+ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and3_1
Xfanout632 _04779_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout643 _03834_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12488__A1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout954_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_4
Xfanout665 net667 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__buf_2
Xfanout676 net677 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout687 net688 vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__buf_2
X_09848_ _04611_ _04670_ _04784_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11160__B2 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\]
+ net957 vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11810_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net270 net267 vssd1 vssd1 vccd1
+ vccd1 _07292_ sky130_fd_sc_hd__a21o_1
XANTENNA__15106__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12790_ _07518_ _07666_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__or2_4
XANTENNA__14010__A _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11741_ _06784_ _07229_ _07198_ _07227_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_1_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11463__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14945__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10671__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14460_ net1278 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__inv_2
X_11672_ net572 _06794_ _07160_ _06271_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_138_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13411_ _07744_ _07836_ _07831_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__o21ba_1
X_10623_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__or4bb_1
XANTENNA__11640__Y _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17293__1349 vssd1 vssd1 vccd1 vccd1 _17293__1349/HI net1349 sky130_fd_sc_hd__conb_1
XFILLER_0_165_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12412__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14391_ net1471 vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_76_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13060__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ _07766_ _07767_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16130_ clknet_leaf_145_wb_clk_i _01799_ _00359_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input83_A wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06108_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11620__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08154__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ net94 team_04_WB.ADDR_START_VAL_REG\[3\] net977 vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__mux2_1
X_16061_ clknet_leaf_129_wb_clk_i _01730_ _00290_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ _06050_ _06060_ _06057_ _06051_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ net1189 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__inv_2
X_12224_ net1967 net510 _07553_ net460 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a22o_1
XANTENNA__12715__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10726__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__X _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ net229 net2475 net513 vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__mux2_1
X_11106_ net531 _06242_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nand2_1
X_16963_ clknet_leaf_125_wb_clk_i _02632_ _01192_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\]
+ sky130_fd_sc_hd__dfrtp_1
X_12086_ net245 net677 vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__and2_1
XANTENNA__12479__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15914_ clknet_leaf_38_wb_clk_i _01591_ _00141_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13140__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ net645 net581 _06252_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11687__C1 _07016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16894_ clknet_leaf_129_wb_clk_i _02563_ _01123_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11151__A1 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15845_ clknet_leaf_87_wb_clk_i _01522_ _00072_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15776_ net1285 vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08329__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ _07640_ _07668_ net317 net1877 vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ net1143 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__inv_2
X_11939_ net1937 net528 net453 _07403_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a22o_1
XANTENNA__12651__A1 _07622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11831__X _07310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09949__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14658_ net1255 vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__inv_2
XANTENNA__08853__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] net1102 vssd1
+ vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__nor2_1
XANTENNA__10594__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12403__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14589_ net1178 vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08702__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__A1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16328_ clknet_leaf_118_wb_clk_i _01997_ _00557_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12094__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16259_ clknet_leaf_117_wb_clk_i _01928_ _00488_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput202 net202 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_11_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12706__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10193__A2 _05800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\]
+ net933 vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13131__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\]
+ net970 vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__mux2_1
X_07894_ team_04_WB.ADDR_START_VAL_REG\[30\] vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__inv_2
XANTENNA__09886__A2 _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__C1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07932__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__mux2_1
XANTENNA__09850__C _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15922__Q net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout368_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09564_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_8__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08515_ net727 _04125_ net712 vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_110_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09495_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10653__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ net751 net717 _03726_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11850__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08377_ net779 _03987_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout702_A net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout323_X net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12158__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10270_ _05865_ _05866_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10533__A team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout440 net443 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 net452 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__clkbuf_4
Xfanout462 _06204_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_4
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_4
X_13960_ net154 net1064 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__and2_1
Xfanout484 net485 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__buf_8
XANTENNA__09533__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _07613_ net328 net384 net1762 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a22o_1
X_13891_ _03195_ _03269_ _03169_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10341__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15630_ net1197 vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__inv_2
X_12842_ _07540_ net346 net395 net1878 vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__a22o_1
XANTENNA__12179__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15561_ net1134 vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__inv_2
XANTENNA__12633__A1 _07604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773_ _07500_ net338 net396 net1635 vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a22o_1
XANTENNA__14675__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17300_ net1356 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
X_14512_ net1191 vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08932__S0 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11724_ _07198_ _07201_ _07202_ _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__and4bb_1
XANTENNA__09769__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15492_ net1171 vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17231_ net1437 _02841_ _01489_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_14443_ net1277 vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__inv_2
X_11655_ _06589_ _07143_ net586 vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12195__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249__1309 vssd1 vssd1 vccd1 vccd1 _17249__1309/HI net1309 sky130_fd_sc_hd__conb_1
XFILLER_0_138_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10606_ net67 net66 _06141_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__or4_1
X_17162_ clknet_leaf_85_wb_clk_i _02774_ _01391_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_88_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12936__A2 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14374_ net1489 vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__clkbuf_1
X_11586_ net465 _07073_ _07074_ _06205_ _07072_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16113_ clknet_leaf_175_wb_clk_i _01782_ _00342_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13325_ team_04_WB.MEM_SIZE_REG_REG\[17\] _07749_ _07750_ vssd1 vssd1 vccd1 vccd1
+ _07751_ sky130_fd_sc_hd__a21o_1
X_10537_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[21\]
+ _06096_ net1049 vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17093_ clknet_leaf_91_wb_clk_i _02728_ _01322_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12149__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09708__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16044_ clknet_leaf_107_wb_clk_i _01713_ _00273_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10468_ _06020_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__nand2_1
X_13256_ net81 team_04_WB.ADDR_START_VAL_REG\[20\] net975 vssd1 vssd1 vccd1 vccd1
+ _01650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10714__Y _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12207_ net249 net650 vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__and2_1
X_13187_ _07623_ net383 net293 net1695 vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a22o_1
XANTENNA__12134__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10399_ _05526_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12138_ net246 net2496 net511 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13113__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16946_ clknet_leaf_8_wb_clk_i _02615_ _01175_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\]
+ sky130_fd_sc_hd__dfrtp_1
X_12069_ net2133 net353 _07489_ net445 vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10332__C1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16877_ clknet_leaf_42_wb_clk_i _02546_ _01106_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\]
+ sky130_fd_sc_hd__dfrtp_1
X_15828_ clknet_leaf_92_wb_clk_i _01505_ _00055_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15759_ net1290 vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__inv_2
XANTENNA__14585__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08300_ _03907_ _03908_ _03909_ _03910_ net828 net735 vssd1 vssd1 vccd1 vccd1 _03911_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09280_ _04885_ _04890_ net771 vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08583__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08231_ net725 _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_74 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12388__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08056__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08162_ net771 _03772_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14129__B2 team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__mux2_1
XANTENNA__12392__X _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11__f_wb_clk_i_X clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xclkload50 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_8
XFILLER_0_141_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload61 clknet_leaf_39_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_77_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09005__B1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload72 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload72/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__13888__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload83 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload83/Y sky130_fd_sc_hd__inv_6
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload94 clknet_leaf_148_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__inv_6
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12560__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__mux2_1
XANTENNA__09308__A1 net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout485_A net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_10_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17292__1348 vssd1 vssd1 vccd1 vccd1 _17292__1348/HI net1348 sky130_fd_sc_hd__conb_1
XANTENNA__14112__X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ net1010 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_3_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09353__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07877_ net1191 vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__inv_2
XANTENNA__08110__X _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout273_X net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10874__B1 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\]
+ net890 vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11418__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\]
+ net951 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout917_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08295__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__mux2_1
XANTENNA__12091__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08429_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12446__C net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload0 clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__12918__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11440_ net574 net561 _05475_ _06208_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__a41o_1
XFILLER_0_163_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11371_ _06512_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ net619 _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nor2_1
X_13110_ _07542_ net370 net298 net1636 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22o_1
X_14090_ net1462 _06126_ net1034 vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__mux2_1
XANTENNA__13558__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _07502_ net382 net309 net1768 vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a22o_1
X_10253_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _05537_ vssd1
+ vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__xor2_1
XANTENNA_input46_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _05542_ vssd1
+ vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__xor2_2
Xfanout1202 net1254 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__clkbuf_2
Xfanout1213 net1220 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
Xfanout1224 net1253 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__buf_2
X_16800_ clknet_leaf_138_wb_clk_i _02469_ _01029_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1235 net1243 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13574__A team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1246 net1252 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1257 net1297 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_4
X_14992_ net1163 vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_135_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout270 _07237_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__clkbuf_2
Xfanout1268 net1280 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout281 _05523_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout1279 net1280 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__buf_2
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_8
X_16731_ clknet_leaf_100_wb_clk_i _02400_ _00960_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\]
+ sky130_fd_sc_hd__dfrtp_1
X_13943_ _03079_ _03080_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or2_1
XANTENNA__10314__C1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ clknet_leaf_14_wb_clk_i _02331_ _00891_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\]
+ sky130_fd_sc_hd__dfrtp_1
X_13874_ _03254_ _03257_ net1834 net1068 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a2bb2o_1
X_15613_ net1154 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__inv_2
X_12825_ _07523_ net340 net394 net1697 vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a22o_1
XANTENNA_output202_A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16593_ clknet_leaf_180_wb_clk_i _02262_ _00822_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15544_ net1205 vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__inv_2
X_12756_ _07481_ net349 net403 net2454 vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7__f_wb_clk_i_X clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_155_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ net464 _07186_ _07195_ net287 vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__a22o_2
XANTENNA__12129__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15475_ net1234 vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ net701 _06183_ _07663_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__or3_4
XFILLER_0_155_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17214_ net1420 _02824_ _01455_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09665__A1_N net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ net1289 vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__inv_2
XANTENNA__08038__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12909__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11638_ _06268_ _06789_ _07124_ _06277_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17145_ clknet_leaf_81_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[1\]
+ _01374_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14357_ net1258 vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__inv_2
Xwire660 _03948_ vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_2
X_11569_ net754 _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__and2_1
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold707 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\] vssd1 vssd1
+ vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ team_04_WB.MEM_SIZE_REG_REG\[25\] _07732_ _07733_ vssd1 vssd1 vccd1 vccd1
+ _07734_ sky130_fd_sc_hd__a21o_1
Xhold718 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\] vssd1 vssd1
+ vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ clknet_leaf_45_wb_clk_i _00024_ _01305_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold729 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\] vssd1 vssd1
+ vccd1 vccd1 net2166 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08342__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14288_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\] _03457_
+ net821 vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_55_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11269__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ clknet_leaf_92_wb_clk_i _01696_ _00256_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13239_ net91 team_04_WB.MEM_SIZE_REG_REG\[2\] net985 vssd1 vssd1 vccd1 vccd1 _01664_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11345__A1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12799__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08780_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16929_ clknet_leaf_133_wb_clk_i _02598_ _01158_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09401_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__mux2_1
XANTENNA__09149__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09332_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12073__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09202__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ net771 _04873_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__nor2_1
XANTENNA__10348__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A2 _07182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08214_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
XANTENNA__09696__X _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08145_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14107__X net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout400_A _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12781__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload150 clknet_leaf_77_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload150/Y sky130_fd_sc_hd__inv_6
X_08076_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__mux2_1
Xclkload161 clknet_leaf_104_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload161/X sky130_fd_sc_hd__clkbuf_4
Xclkload172 clknet_leaf_85_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload172/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12282__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__C1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09529__A1 _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11336__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_164_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 net138 vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\] vssd1 vssd1 vccd1
+ vccd1 net1471 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08488__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__mux2_1
Xhold45 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[9\]
+ vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09083__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248__1308 vssd1 vssd1 vccd1 vccd1 _17248__1308/HI net1308 sky130_fd_sc_hd__conb_1
Xhold56 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\] vssd1 vssd1 vccd1
+ vccd1 net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[7\] vssd1 vssd1
+ vccd1 vccd1 net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[5\] vssd1
+ vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\] _03524_
+ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__nor2_1
XANTENNA__10530__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 net124 vssd1 vssd1 vccd1 vccd1 net1526 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout655_X net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08060__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _04865_ _04919_ _04973_ _06286_ net659 vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__a41o_1
XFILLER_0_98_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10311__A2 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10871_ _04585_ _06358_ _06359_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__nand3_1
XFILLER_0_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input100_A wbs_dat_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _07579_ net482 net412 net1896 vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a22o_1
XANTENNA__13261__A1 team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ _02971_ _02975_ _02978_ team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1
+ vccd1 _02981_ sky130_fd_sc_hd__a31o_1
XANTENNA__08427__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ net2131 net243 net420 vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11811__A2 _07292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13013__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15260_ net1148 vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12472_ net525 net611 _07473_ net431 net1825 vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ net1088 net1087 _03406_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__a31o_1
X_11423_ net568 _06716_ _06251_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__a21o_1
X_15191_ net1230 vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] _03363_
+ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__nor2_1
X_11354_ _06348_ _06354_ _06657_ net463 vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10705__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10305_ net623 _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14073_ net1486 _06092_ net1032 vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__mux2_1
X_11285_ net564 _06246_ _06612_ _06271_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ net280 _05835_ _05838_ _05525_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__o22a_1
X_13024_ _07485_ net373 net307 net1638 vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a22o_1
Xfanout1010 _03547_ vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_2
Xfanout1021 _06073_ vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__clkbuf_2
Xfanout1032 net1035 vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_4
X_10167_ net622 _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__nor2_1
Xfanout1043 net1044 vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__buf_2
Xfanout1054 _03541_ vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_2
Xfanout1065 _07700_ vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_2
Xfanout1076 _03525_ vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__buf_4
Xfanout1087 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_2
X_10098_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _04786_ vssd1
+ vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__or2_1
X_14975_ net1266 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__inv_2
Xfanout1098 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\] vssd1
+ vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_2
XFILLER_0_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16714_ clknet_leaf_161_wb_clk_i _02383_ _00943_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\]
+ sky130_fd_sc_hd__dfrtp_1
X_13926_ net1662 net1071 _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10302__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09721__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16645_ clknet_leaf_4_wb_clk_i _02314_ _00874_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\]
+ sky130_fd_sc_hd__dfrtp_1
X_13857_ net1663 net1066 _03231_ _03246_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12808_ net256 net2576 net325 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__mux2_1
X_16576_ clknet_leaf_139_wb_clk_i _02245_ _00805_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13788_ team_04_WB.ADDR_START_VAL_REG\[17\] _03171_ _03175_ _03178_ vssd1 vssd1 vccd1
+ vccd1 _03179_ sky130_fd_sc_hd__and4_1
X_15527_ net1141 vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__inv_2
XANTENNA__11263__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _07464_ net348 net403 net2505 vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_32_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09957__A _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15458_ net1240 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__inv_2
XANTENNA__13004__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17291__1347 vssd1 vssd1 vccd1 vccd1 _17291__1347/HI net1347 sky130_fd_sc_hd__conb_1
XFILLER_0_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ net1267 vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14074__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15389_ net1153 vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__inv_2
XANTENNA__12763__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17128_ clknet_leaf_76_wb_clk_i net1509 _01357_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold504 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\] vssd1 vssd1
+ vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08072__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold515 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\] vssd1 vssd1
+ vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold526 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\] vssd1 vssd1
+ vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\] vssd1 vssd1
+ vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold548 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\] vssd1 vssd1
+ vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ clknet_leaf_48_wb_clk_i _00037_ _01288_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_09950_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__inv_2
Xhold559 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\] vssd1 vssd1
+ vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09606__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08901_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ net590 net633 vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_70_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11727__A net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\] _03650_ _03652_
+ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1204 _00031_ vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1215 team_04_WB.instance_to_wrap.final_design.uart.receiving vssd1 vssd1 vccd1
+ vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1226 team_04_WB.ADDR_START_VAL_REG\[30\] vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08763_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13491__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08694_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\]
+ net941 vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XANTENNA__13491__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09631__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__A_N net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12046__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__mux2_1
XANTENNA__13794__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout615_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10509__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07939__X _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ _04853_ _04854_ _04855_ _04856_ net826 net734 vssd1 vssd1 vccd1 vccd1 _04857_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08128_ _03735_ _03736_ _03737_ _03738_ net825 net733 vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12754__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout984_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__mux2_1
XANTENNA__12506__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09806__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _03946_ net549 _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 wbs_we_i vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
X_10021_ _05585_ _05631_ _05586_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16001__Q team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14760_ net1124 vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__inv_2
XANTENNA__08489__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15784__3 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__inv_2
X_11972_ net695 _07089_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12285__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08946__A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13711_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] net1045 _03101_
+ _03515_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__o22a_1
X_10923_ _06410_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14691_ net1172 vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13063__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16430_ clknet_leaf_27_wb_clk_i _02099_ _00659_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13642_ _07794_ _07795_ _07797_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__o21ba_1
XANTENNA__09113__Y _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__inv_2
XANTENNA__12187__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11245__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16361_ clknet_leaf_100_wb_clk_i _02030_ _00590_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\]
+ sky130_fd_sc_hd__dfrtp_1
X_13573_ _02961_ _02963_ net998 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ net561 _06245_ _06263_ _06266_ _06273_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__o221a_1
XANTENNA__11796__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12993__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15312_ net1162 vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ net2119 net214 net422 vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16292_ clknet_leaf_167_wb_clk_i _01961_ _00521_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13299__A _06592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15243_ net1161 vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__inv_2
X_12455_ net2390 net428 _07647_ net520 vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a22o_1
XANTENNA__10716__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12745__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11406_ net534 _06894_ _06893_ net564 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_10_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15174_ net1104 vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12386_ net223 net2432 net497 vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10220__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14125_ team_04_WB.MEM_SIZE_REG_REG\[24\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[24\]
+ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__a22o_1
XFILLER_0_132_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _06791_ _06797_ net554 vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_150_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_150_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_91_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09716__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ net31 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1
+ vccd1 vccd1 _01530_ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11268_ _06734_ net284 vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__nor2_1
XANTENNA__13170__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13238__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ net611 _07467_ net474 net313 net1783 vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a32o_1
X_10219_ _05540_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__nor2_1
XANTENNA__12142__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08272__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ _06485_ _06687_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14958_ net1197 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09451__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ net1042 _03282_ _03283_ net1067 net1517 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a32o_1
XANTENNA__10597__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14889_ net1133 vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_46_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11282__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16628_ clknet_leaf_2_wb_clk_i _02297_ _00857_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13225__A1 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12028__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15689__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09524__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16559_ clknet_leaf_189_wb_clk_i _02228_ _00788_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ net780 _04710_ net763 vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__o21a_1
XANTENNA__12984__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09031_ _04612_ _04641_ net666 vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux2_2
X_17247__1307 vssd1 vssd1 vccd1 vccd1 _17247__1307/HI net1307 sky130_fd_sc_hd__conb_1
XFILLER_0_150_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11539__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold301 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\] vssd1 vssd1
+ vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12200__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold312 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\] vssd1 vssd1
+ vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\] vssd1 vssd1
+ vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\] vssd1 vssd1
+ vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold345 net121 vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold356 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\] vssd1 vssd1
+ vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold367 team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09626__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold378 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\] vssd1 vssd1
+ vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] _05543_ vssd1
+ vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__xor2_2
Xhold389 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\] vssd1 vssd1
+ vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout803 _03551_ vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__buf_4
XANTENNA__15925__Q net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout814 net815 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
Xfanout825 net830 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout836 net837 vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_4
Xfanout847 net859 vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
X_09864_ _05378_ net532 vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__nor2_2
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_2
Xfanout869 net870 vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_4
Xhold1001 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\] vssd1 vssd1
+ vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\] vssd1 vssd1
+ vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ net776 _04419_ net764 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__o21a_1
Xhold1023 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\] vssd1 vssd1
+ vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[8\] team_04_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ net1010 vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__mux2_1
Xhold1034 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\] vssd1 vssd1
+ vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\] vssd1 vssd1
+ vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\] vssd1 vssd1
+ vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14110__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1067 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\] vssd1 vssd1
+ vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ net661 _04355_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__o21ai_4
Xhold1078 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\] vssd1 vssd1
+ vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12267__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08766__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\] vssd1 vssd1
+ vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13391__B team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__B1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08677_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout353_X net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1095_X net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08891__A1 _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout520_X net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_X net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12975__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10570_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[10\]
+ _06118_ net1048 vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08705__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09229_ net666 _04839_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__nor2_1
XANTENNA__12990__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10536__A team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14008__A _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12727__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__C net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ net226 net672 vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12171_ net227 net648 vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11122_ net584 _06610_ net289 vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__o21a_1
XANTENNA__08440__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold890 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\] vssd1 vssd1
+ vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13058__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15930_ clknet_leaf_59_wb_clk_i _01607_ _00157_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfrtp_1
X_11053_ _06540_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__nand2_1
X_10004_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15861_ clknet_leaf_94_wb_clk_i _01538_ _00088_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_17290__1346 vssd1 vssd1 vccd1 vccd1 _17290__1346/HI net1346 sky130_fd_sc_hd__conb_1
X_14812_ net1126 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14743_ net1226 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__inv_2
XANTENNA__11814__B net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11955_ _03631_ _05981_ net696 _07416_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10906_ net580 _06394_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14674_ net1237 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11886_ net757 _05910_ _06185_ _04612_ net690 vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__o221a_1
XANTENNA__11481__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16413_ clknet_leaf_129_wb_clk_i _02082_ _00642_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\]
+ sky130_fd_sc_hd__dfrtp_1
X_13625_ team_04_WB.ADDR_START_VAL_REG\[6\] _03014_ vssd1 vssd1 vccd1 vccd1 _03016_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13758__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10837_ _03891_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12966__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16344_ clknet_leaf_153_wb_clk_i _02013_ _00573_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13556_ _02909_ _02945_ _02946_ _02922_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_41_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08634__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _05449_ net467 _05469_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__and3_4
XFILLER_0_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12507_ _07504_ net486 net424 net1976 vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16275_ clknet_leaf_184_wb_clk_i _01944_ _00504_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12137__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ _07864_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__xor2_1
XANTENNA__12981__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10699_ _03621_ net691 vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__nor2_1
XANTENNA__12718__B1 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15226_ net1138 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12438_ net611 _07446_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_130_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12194__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15157_ net1207 vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ net247 net2464 net495 vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11941__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14108_ team_04_WB.MEM_SIZE_REG_REG\[7\] net988 net981 team_04_WB.ADDR_START_VAL_REG\[7\]
+ net1005 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__o221a_2
XTAP_TAPCELL_ROW_39_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15088_ net1163 vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13143__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ net18 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1
+ vccd1 vccd1 _01547_ sky130_fd_sc_hd__a22o_1
XANTENNA__12497__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08600_ _04207_ _04208_ _04209_ _04210_ net783 net805 vssd1 vssd1 vccd1 vccd1 _04211_
+ sky130_fd_sc_hd__mux4_1
X_09580_ net718 _05190_ _05179_ _05178_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__12249__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08531_ net594 _04139_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08548__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13997__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_100_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08462_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ net751 _04002_ _03725_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_102_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10680__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_169_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12957__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_154_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07979__A3 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout313_A _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1055_A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12709__B1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10075__B _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold120 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1557 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13667__A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold131 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\] vssd1 vssd1
+ vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\] vssd1 vssd1
+ vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\] vssd1 vssd1
+ vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09356__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\] vssd1 vssd1
+ vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08113__X _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\] vssd1 vssd1
+ vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[27\] vssd1
+ vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12290__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\] vssd1 vssd1
+ vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net602 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__buf_2
XANTENNA__13134__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
X_09916_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05526_ vssd1
+ vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__and2_1
Xfanout622 net624 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_2
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout633 _04779_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08236__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12488__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__buf_4
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__buf_4
X_09847_ _05455_ _05457_ _03621_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__o21a_1
Xfanout677 _07482_ vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_4
Xfanout688 _06199_ vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_2
XANTENNA_fanout470_X net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14498__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__mux2_1
XANTENNA__09091__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11740_ _06709_ _06710_ _06761_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_1_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_189_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10671__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _07157_ _07159_ net572 vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12948__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ net1084 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 _07836_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10622_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\]
+ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08435__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14390_ net1461 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12412__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] team_04_WB.MEM_SIZE_REG_REG\[11\]
+ _07765_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ _06107_ net1637 net1021 vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
XANTENNA__12963__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16060_ clknet_leaf_129_wb_clk_i _01729_ _00289_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_13272_ net95 team_04_WB.ADDR_START_VAL_REG\[4\] net977 vssd1 vssd1 vccd1 vccd1 _01634_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input76_A wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10484_ _06013_ _06047_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_161_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15011_ net1175 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__inv_2
XANTENNA__12176__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _07443_ _07444_ net650 vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11923__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ net231 net2602 net513 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
XANTENNA__08023__X _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13125__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _06237_ _06244_ net537 vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__mux2_1
X_12085_ net2182 net353 _07497_ net447 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a22o_1
X_16962_ clknet_leaf_147_wb_clk_i _02631_ _01191_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12479__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _06493_ _06524_ net464 vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__o21ai_1
X_15913_ clknet_leaf_124_wb_clk_i _01590_ _00140_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16893_ clknet_leaf_132_wb_clk_i _02562_ _01122_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15844_ clknet_leaf_88_wb_clk_i _01521_ _00071_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_17246__1306 vssd1 vssd1 vccd1 vccd1 _17246__1306/HI net1306 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_86_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15775_ net1288 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__inv_2
XANTENNA__13979__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ _07639_ net474 net316 net1936 vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14726_ net1104 vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ net653 net261 vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__and2_2
XANTENNA__12651__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10662__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14657_ net1148 vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11869_ net705 _05892_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_60_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12939__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13251__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13608_ _07024_ net271 _07687_ _02998_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14588_ net1184 vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__inv_2
XANTENNA__12403__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08345__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10414__A1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16327_ clknet_leaf_164_wb_clk_i _01996_ _00556_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13539_ team_04_WB.ADDR_START_VAL_REG\[21\] _02923_ _02929_ vssd1 vssd1 vccd1 vccd1
+ _02930_ sky130_fd_sc_hd__and3_1
XANTENNA__08702__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09965__A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16258_ clknet_leaf_143_wb_clk_i _01927_ _00487_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput203 net203 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
X_15209_ net1135 vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__inv_2
XANTENNA__14082__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ clknet_leaf_141_wb_clk_i _01858_ _00418_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11914__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13116__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07962_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ net625 net555 vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_147_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07893_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\] vssd1 vssd1
+ vccd1 vccd1 _03508_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_74_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07932__B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__D net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09718__S0 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout263_A _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08514_ _04121_ _04122_ _04123_ _04124_ net824 net733 vssd1 vssd1 vccd1 vccd1 _04125_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_19_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09494_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\]
+ net949 vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__mux2_1
XANTENNA__12642__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10653__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08445_ net751 net717 _03726_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout430_A _07641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1172_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout528_A _06195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08376_ _03983_ _03984_ _03985_ _03986_ net784 net805 vssd1 vssd1 vccd1 vccd1 _03987_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13949__X _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14781__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07947__X _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09875__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08457__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout430 _07641_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_4
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__clkbuf_4
Xfanout452 net461 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
Xfanout463 _06204_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_92_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout474 _07668_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_4
Xfanout485 net486 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout496 _07624_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_6
X_12910_ _07612_ net337 net384 net1931 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__a22o_1
XANTENNA__12330__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ _03148_ _03193_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__or2_1
XANTENNA__12881__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ _07539_ net348 net395 net2162 vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ net1116 vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__inv_2
X_12772_ _07499_ net346 net399 net2636 vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
XANTENNA__12633__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14511_ net1259 vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11723_ _06684_ _07205_ _07211_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__nor3_1
XFILLER_0_138_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11841__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15491_ net1170 vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__inv_2
XANTENNA__08932__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13071__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17230_ net1436 _02840_ _01487_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_83_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ net1272 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__inv_2
XANTENNA__08165__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ net574 _06666_ _07142_ _06250_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__o211a_1
XFILLER_0_166_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12195__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ net65 net64 net47 net36 vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__or4_1
XANTENNA__13594__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17161_ clknet_leaf_85_wb_clk_i _02773_ _01390_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12397__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14373_ net1474 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11585_ _06395_ _06422_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__or2_1
X_16112_ clknet_leaf_0_wb_clk_i _01781_ _00341_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13324_ _07747_ _07748_ _07749_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__o21ba_1
X_17092_ clknet_leaf_43_wb_clk_i _02727_ _01321_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10536_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] net1097 net1053 vssd1 vssd1 vccd1
+ vccd1 _06096_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output182_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16043_ clknet_leaf_22_wb_clk_i _01712_ _00272_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_13255_ net82 team_04_WB.ADDR_START_VAL_REG\[21\] net975 vssd1 vssd1 vccd1 vccd1
+ _01651_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ _06028_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12206_ net2226 net507 _07544_ net441 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_36_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13186_ _07622_ net380 net292 net1712 vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a22o_1
X_10398_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\]
+ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] vssd1 vssd1 vccd1 vccd1
+ _05982_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_36_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12137_ net236 net2442 net511 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08688__X _04299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__S net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16945_ clknet_leaf_179_wb_clk_i _02614_ _01174_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\]
+ sky130_fd_sc_hd__dfrtp_1
X_12068_ net217 net677 vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11019_ team_04_WB.MEM_SIZE_REG_REG\[15\] team_04_WB.MEM_SIZE_REG_REG\[14\] _06507_
+ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__or3_1
XANTENNA__15027__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12003__X _07455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16876_ clknet_leaf_120_wb_clk_i _02545_ _01105_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12872__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15827_ clknet_leaf_91_wb_clk_i _01504_ _00054_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__X _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15758_ net1283 vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__inv_2
XANTENNA__08828__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12624__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ net1199 vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__inv_2
XANTENNA__14077__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15689_ net1257 vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08230_ _03837_ _03838_ _03839_ _03840_ net831 net737 vssd1 vssd1 vccd1 vccd1 _03841_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _03768_ _03769_ _03770_ _03771_ net786 net807 vssd1 vssd1 vccd1 vccd1 _03772_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09253__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11596__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14129__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ net771 _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload40 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload51 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__clkinv_4
Xclkload62 clknet_leaf_43_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload62/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload73 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload73/X sky130_fd_sc_hd__clkbuf_8
Xclkload84 clknet_leaf_57_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_6
Xclkload95 clknet_leaf_149_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload95/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11899__B1 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_149_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08994_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__mux2_1
XANTENNA__09634__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09308__A2 _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] net1010 vssd1 vssd1 vccd1 vccd1
+ _03556_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12863__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09615_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__mux2_1
XANTENNA__12615__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11912__B _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09477_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\]
+ net947 vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout812_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_X net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13576__B1 team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload1 clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__inv_8
XFILLER_0_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__mux2_1
XANTENNA__13040__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11051__A1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ team_04_WB.MEM_SIZE_REG_REG\[20\] _06511_ team_04_WB.MEM_SIZE_REG_REG\[21\]
+ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08713__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17245__1305 vssd1 vssd1 vccd1 vccd1 _17245__1305/HI net1305 sky130_fd_sc_hd__conb_1
XFILLER_0_6_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ _05631_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14016__A _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13040_ _07501_ net383 net308 net2201 vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a22o_1
X_10252_ net620 _05848_ _05852_ net280 vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12551__A1 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16004__Q team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _05787_ _05788_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__o21ai_1
Xfanout1203 net1206 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 net1216 vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__buf_4
XANTENNA__09544__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1225 net1227 vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__buf_4
Xfanout1236 net1243 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input39_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ net1140 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__inv_2
Xfanout1247 net1252 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_2
Xfanout1258 net1261 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 _07327_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__clkbuf_2
Xfanout271 _07216_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_4
Xfanout1269 net1280 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__buf_2
XANTENNA__13066__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout282 _05523_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_4
X_13942_ _03083_ net1041 _03303_ net1073 net1529 vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__a32o_1
X_16730_ clknet_leaf_37_wb_clk_i _02399_ _00959_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout293 _07684_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08020__Y _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ clknet_leaf_33_wb_clk_i _02330_ _00890_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\]
+ sky130_fd_sc_hd__dfrtp_1
X_13873_ _03200_ _03220_ net1039 vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_175_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_175_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14056__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15612_ net1147 vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12824_ _07522_ net334 net393 net1884 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a22o_1
XANTENNA__12067__B1 _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16592_ clknet_leaf_191_wb_clk_i _02261_ _00821_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12606__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15543_ net1233 vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12755_ _07480_ net345 net402 net2189 vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11706_ _07187_ _07193_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__and3_1
X_15474_ net1247 vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12686_ _05111_ _06189_ _06191_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__or3b_4
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17213_ net1419 _02823_ _01453_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_14425_ net1283 vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__inv_2
X_11637_ _05110_ net587 net359 _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_154_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08669__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17144_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[0\]
+ _01373_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09719__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ net1258 vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11568_ _07042_ _07055_ _07056_ _07041_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__a31oi_4
XANTENNA__08623__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ _07730_ _07731_ _07732_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold708 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\] vssd1 vssd1
+ vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
X_17075_ clknet_leaf_45_wb_clk_i _00023_ _01304_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10519_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[27\]
+ _06084_ net1048 vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__mux2_1
Xhold719 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\] vssd1 vssd1
+ vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
X_14287_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\] _03457_
+ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__and2_1
XANTENNA__12145__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ net569 _06768_ _06251_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_139_Left_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16026_ clknet_leaf_77_wb_clk_i _00002_ _00255_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_55_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13238_ net94 team_04_WB.MEM_SIZE_REG_REG\[3\] net984 vssd1 vssd1 vccd1 vccd1 _01665_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11984__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10604__D net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _07605_ net373 net291 net1947 vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__a22o_1
XANTENNA__08859__A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__X _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16928_ clknet_leaf_138_wb_clk_i _02597_ _01157_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12845__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16859_ clknet_leaf_97_wb_clk_i _02528_ _01088_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14047__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Left_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09400_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__mux2_1
XANTENNA__09149__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08594__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[552\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09262_ _04869_ _04870_ _04871_ _04872_ net786 net807 vssd1 vssd1 vccd1 vccd1 _04873_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08213_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09193_ _04800_ _04801_ _04802_ _04803_ net826 net734 vssd1 vssd1 vccd1 vccd1 _04804_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13022__A2 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout226_A _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15220__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09629__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _03696_ _03754_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nand2_1
XANTENNA__08533__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_157_Left_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload140 clknet_leaf_119_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload140/Y sky130_fd_sc_hd__inv_8
X_08075_ _03682_ _03683_ _03684_ _03685_ net827 net735 vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload151 clknet_leaf_79_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload151/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1135_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload162 clknet_leaf_120_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload162/Y sky130_fd_sc_hd__clkinv_2
Xclkload173 clknet_leaf_86_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload173/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_168_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09529__A2 _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12533__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout595_A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07944__Y _03555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14123__X net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold13 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\] vssd1 vssd1 vccd1
+ vccd1 net1450 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\] vssd1 vssd1 vccd1
+ vccd1 net1461 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout762_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\] vssd1 vssd1
+ vccd1 vccd1 net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11195__A _06681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold57 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[7\]
+ vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ net1077 net1031 vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_1
Xhold68 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _02765_ vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12836__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10530__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_166_Left_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09725__A1_N net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14038__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ _04642_ _05463_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08708__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _03634_ _05137_ _05138_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15801__20 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__inv_2
XANTENNA__10539__A team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ net2211 net255 net423 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12471_ net520 net602 _07472_ net428 net1940 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14210_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__inv_2
XFILLER_0_151_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09539__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ _06870_ _06910_ net561 vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__mux2_1
XANTENNA__08443__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15190_ net1224 vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__inv_2
X_14141_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[8\]
+ _03522_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11353_ _06348_ _06657_ _06354_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10304_ _05755_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__xnor2_1
X_14072_ net1514 _06090_ net1034 vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11284_ net568 _06698_ _06772_ net583 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__a211o_1
XANTENNA__12524__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13023_ net699 _07483_ _07666_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__or3_4
X_10235_ net1055 _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__nor2_1
Xfanout1000 _07686_ vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__clkbuf_2
Xfanout1011 _03547_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_4
Xfanout1022 _06073_ vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__clkbuf_4
Xfanout1033 net1035 vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
X_10166_ _05775_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__xnor2_1
Xfanout1044 net1046 vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__buf_2
Xfanout1055 net1056 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__clkbuf_4
Xfanout1066 net1067 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_2
Xfanout1077 _03524_ vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1088 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_2
X_10097_ _05706_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12827__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14974_ net1239 vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__inv_2
Xfanout1099 net1100 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__clkbuf_4
X_16713_ clknet_leaf_122_wb_clk_i _02382_ _00942_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\]
+ sky130_fd_sc_hd__dfrtp_1
X_13925_ _03132_ _03140_ _03292_ net1040 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__o31a_1
XFILLER_0_156_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload4_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ _02855_ _03228_ _03230_ _03243_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a31oi_1
X_16644_ clknet_leaf_171_wb_clk_i _02313_ _00873_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12807_ net258 net2544 net324 vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
XANTENNA__11552__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13787_ net998 _03177_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__nand2_1
X_16575_ clknet_leaf_157_wb_clk_i _02244_ _00804_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10999_ _06327_ _06330_ _06332_ _06484_ _06326_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__a221o_1
XANTENNA__11799__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11263__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12738_ _07463_ net334 net401 net2360 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a22o_1
X_15526_ net1103 vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__inv_2
XANTENNA__12460__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12935__Y _07676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15457_ net1130 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ net259 net2278 net476 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14408_ net1277 vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09449__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15040__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_72_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_160_Right_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ net1145 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__inv_2
XANTENNA__08353__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_17127_ clknet_leaf_76_wb_clk_i net1522 _01356_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14339_ net1183 vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold505 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\] vssd1 vssd1
+ vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\] vssd1 vssd1
+ vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\] vssd1 vssd1
+ vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\] vssd1 vssd1
+ vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ clknet_leaf_48_wb_clk_i _00036_ _01287_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold549 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\] vssd1 vssd1
+ vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16009_ clknet_4_5__leaf_wb_clk_i _01685_ _00238_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_08900_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14090__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _04814_ _04865_ net631 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_70_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__or3_1
Xhold1205 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\] vssd1 vssd1
+ vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\] vssd1 vssd1
+ vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1227 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] vssd1 vssd1
+ vccd1 vccd1 net2664 sky130_fd_sc_hd__dlygate4sd3_1
X_08762_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08693_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\]
+ net941 vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17244__1304 vssd1 vssd1 vccd1 vccd1 _17244__1304/HI net1304 sky130_fd_sc_hd__conb_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout343_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09314_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12451__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09245_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout510_A _07521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14118__X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout608_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_X net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09176_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\]
+ net852 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1040_X net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08058_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout977_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _05587_ _05588_ _05628_ _04671_ net634 vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__o32ai_4
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07933__B2 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11971_ net692 _07428_ _07430_ net616 vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_95_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13710_ _07806_ _03100_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__xnor2_1
X_10922_ _06408_ _06409_ _05404_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14690_ net1255 vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__inv_2
XANTENNA__08438__S net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13641_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__inv_2
X_10853_ _04166_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14964__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16360_ clknet_leaf_118_wb_clk_i _02029_ _00589_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\]
+ sky130_fd_sc_hd__dfrtp_1
X_13572_ net994 _02960_ _02962_ net990 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o2bb2a_1
X_10784_ net569 _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__nor2_2
X_15311_ net1196 vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12523_ net2247 net212 net422 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16291_ clknet_leaf_119_wb_clk_i _01960_ _00520_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15242_ net1107 vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__inv_2
XANTENNA__13299__B net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12454_ net601 net240 net680 vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10716__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ net635 _04724_ _05377_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__mux2_1
XANTENNA__13942__B1 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15173_ net1109 vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__inv_2
X_12385_ net234 net2456 net497 vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14124_ team_04_WB.MEM_SIZE_REG_REG\[23\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[23\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__o221a_1
X_11336_ net582 _06532_ _06824_ net288 vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__o31a_1
XANTENNA__08901__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14055_ net32 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1
+ vccd1 vccd1 _01531_ sky130_fd_sc_hd__a22o_1
XANTENNA__11828__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ _06748_ _06750_ _06755_ _06744_ net286 vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__a2111oi_1
X_13006_ net606 _07466_ net471 net311 net2026 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a32o_1
X_10218_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _05539_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a21oi_1
X_11198_ _06337_ _06482_ _06336_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07924__A1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_190_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_190_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08272__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ _03497_ _04387_ _05759_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__o21bai_1
XANTENNA__13458__C1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11834__Y _07313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14957_ net1152 vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ _02965_ _03281_ _02958_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12681__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14888_ net1116 vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09033__A _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16627_ clknet_leaf_183_wb_clk_i _02296_ _00856_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\]
+ sky130_fd_sc_hd__dfrtp_1
X_13839_ _03222_ _03224_ _03229_ _02900_ _02875_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__o2111ai_2
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11850__X _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09524__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16558_ clknet_leaf_26_wb_clk_i _02227_ _00787_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08872__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15792__11 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11787__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15509_ net1215 vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__inv_2
XANTENNA__12394__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ clknet_leaf_100_wb_clk_i _02158_ _00718_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10907__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09179__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ net719 _04640_ _04629_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_127_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08083__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09288__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11539__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__B1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold302 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\] vssd1 vssd1
+ vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold313 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\] vssd1 vssd1
+ vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10211__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold324 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\] vssd1 vssd1
+ vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[24\]
+ vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08811__S net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\] vssd1 vssd1
+ vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\] vssd1 vssd1
+ vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09932_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\]
+ _05542_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold368 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\] vssd1 vssd1
+ vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\] vssd1 vssd1
+ vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout815 net817 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_2
Xfanout826 net830 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_8
Xfanout837 net838 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
X_09863_ net549 net531 vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nor2_1
XANTENNA__08112__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net859 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_2
XANTENNA__11172__A0 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_A _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net904 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_2
Xhold1002 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\] vssd1 vssd1
+ vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ net781 _04424_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__or2_1
Xhold1013 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\] vssd1 vssd1
+ vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09794_ net759 _03622_ _03635_ _03662_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__o31a_1
Xhold1024 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\] vssd1 vssd1
+ vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\] vssd1 vssd1
+ vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09642__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14110__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1046 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\] vssd1 vssd1
+ vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ net769 net702 _04330_ net663 vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__a211o_1
Xhold1057 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\] vssd1 vssd1
+ vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09668__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1068 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\] vssd1 vssd1
+ vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\] vssd1 vssd1
+ vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12672__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ net727 _04286_ net712 vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12288__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_179_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14784__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12856__X _07673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12424__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12975__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout513_X net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_X net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09089__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _03723_ _03727_ _03630_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09279__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09817__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ net2225 net508 _07526_ net445 vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ net575 _06609_ _06532_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\] vssd1 vssd1
+ vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\] vssd1 vssd1
+ vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11000__X _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _03754_ net364 _06270_ _06530_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o22a_1
XANTENNA__08022__A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _05404_ _05408_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__xor2_1
X_15860_ clknet_leaf_94_wb_clk_i _01537_ _00087_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input21_A DAT_I[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14811_ net1111 vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__inv_2
XANTENNA__15851__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13074__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12663__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ net756 _05983_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__nor2_1
X_14742_ net1225 vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ _05192_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__xnor2_1
X_14673_ net1274 vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net1805 net528 net451 _07357_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_103_Left_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13624_ team_04_WB.ADDR_START_VAL_REG\[6\] _03014_ vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__and2_1
X_16412_ clknet_leaf_116_wb_clk_i _02081_ _00641_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12415__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10836_ _03919_ _06307_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__xor2_1
XANTENNA__13758__A3 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13555_ _02932_ _02941_ _02930_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_15_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16343_ clknet_leaf_166_wb_clk_i _02012_ _00572_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10767_ net645 _03695_ _06255_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_41_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09831__A1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08634__A2 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ _07503_ net491 net426 net2007 vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
X_16274_ clknet_leaf_6_wb_clk_i _01943_ _00503_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _07856_ _07858_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__nand2_1
X_10698_ net759 _03629_ _03635_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16009__CLK clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15225_ net1246 vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__inv_2
X_12437_ net2394 net434 _07639_ net524 vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a22o_1
XANTENNA__10729__A0 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12194__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15156_ net1225 vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__inv_2
XANTENNA__08631__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12368_ net239 net2555 net495 vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14107_ team_04_WB.MEM_SIZE_REG_REG\[6\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[6\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__o221a_2
XANTENNA__13249__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_112_Left_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11319_ net571 _06807_ _06804_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15087_ net1140 vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__inv_2
XANTENNA__12153__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12299_ net215 net670 vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14038_ net19 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1
+ vccd1 vccd1 _01548_ sky130_fd_sc_hd__o22a_1
XANTENNA__13952__A_N _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14869__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15989_ clknet_leaf_78_wb_clk_i _01665_ _00218_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_171_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11293__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ net594 _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nand2_1
XANTENNA__12654__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Left_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08461_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08392_ net751 _04002_ _03725_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_102_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08806__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09013_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_171_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13948__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1547 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[26\] vssd1
+ vssd1 vccd1 vccd1 net1558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08541__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\] vssd1 vssd1
+ vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\] vssd1 vssd1
+ vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11932__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\] vssd1 vssd1
+ vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\] vssd1 vssd1
+ vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[5\]
+ vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1215_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12290__C net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__buf_2
Xhold187 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\] vssd1 vssd1
+ vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\] vssd1 vssd1
+ vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _07251_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__buf_2
X_09915_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\]
+ net1059 vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__and3_1
Xfanout623 net624 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10091__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout634 _04668_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA__13685__A2 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout675_A _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_X net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_4
Xfanout656 _06182_ vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_4
Xfanout667 _03633_ vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_2
X_09846_ _04669_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__nor2_1
XANTENNA__14131__X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout678 net679 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__buf_4
XANTENNA__12893__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout689 net692 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09372__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\]
+ net957 vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__mux2_1
XANTENNA__12645__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11931__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10671__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11670_ net530 _06564_ _07158_ net559 vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10621_ team_04_WB.EN_VAL_REG net69 _06155_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__mux2_1
XANTENNA__10408__C1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__A0 _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] team_04_WB.MEM_SIZE_REG_REG\[11\]
+ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[16\]
+ _06106_ net1048 vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ net96 team_04_WB.ADDR_START_VAL_REG\[5\] net977 vssd1 vssd1 vccd1 vccd1 _01635_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10483_ _06020_ _06055_ _06013_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_129_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15010_ net1265 vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__inv_2
XANTENNA__12176__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ net2195 net509 _07552_ net455 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XANTENNA_input69_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15846__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11923__A2 _06991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13069__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net223 net2525 net513 vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _06490_ _06492_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
X_16961_ clknet_leaf_133_wb_clk_i _02630_ _01190_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\]
+ sky130_fd_sc_hd__dfrtp_1
X_12084_ net260 net677 vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__and2_2
X_11035_ _06318_ _06491_ _06315_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__a21oi_1
X_15912_ clknet_leaf_118_wb_clk_i _01589_ _00139_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12884__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ clknet_leaf_126_wb_clk_i _02561_ _01121_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ clknet_leaf_90_wb_clk_i _01520_ _00070_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_86_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ net1285 vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__inv_2
X_12986_ _07638_ net472 net317 net2075 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a22o_1
XANTENNA__13979__A3 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12636__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14725_ net1113 vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11937_ net691 _07023_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__o21a_4
XFILLER_0_169_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11868_ net757 _05895_ _06185_ _04502_ net690 vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__o221a_1
XANTENNA__10662__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08626__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14656_ net1217 vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09311__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ _07685_ _07691_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_60_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10819_ _03919_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__nor2_1
XANTENNA__12148__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14587_ net1179 vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11799_ net694 _07196_ _07282_ net615 vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10414__A2 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16326_ clknet_leaf_17_wb_clk_i _01995_ _00555_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11072__C1 _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13538_ _02926_ _02928_ net996 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13469_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _05793_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16257_ clknet_leaf_136_wb_clk_i _01926_ _00486_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09568__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09457__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ net1118 vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__inv_2
Xoutput204 net204 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_0_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08361__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16188_ clknet_leaf_128_wb_clk_i _01857_ _00417_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09663__S0 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15139_ net1168 vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07961_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\]
+ net933 vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__mux2_1
X_09700_ net625 net565 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__nand2_1
XANTENNA__12875__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\] vssd1 vssd1
+ vccd1 vccd1 _03507_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08543__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09192__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__mux2_1
X_09562_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12627__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09718__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08513_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\]
+ net846 vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__mux2_1
XANTENNA__13950__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09493_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ net766 _04054_ _04043_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10653__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_173_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13052__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout423_A _07658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout211_X net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08457__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10533__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout420 _07658_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_6
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 _07641_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__buf_2
XANTENNA__13617__S net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10830__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout453 net457 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 _06203_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12866__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout475 _07662_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_6
Xfanout486 net494 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12330__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ _05439_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__inv_2
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_6
XANTENNA__10341__A1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ _07538_ net350 net394 net1704 vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__a22o_1
XANTENNA__12618__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17329__1385 vssd1 vssd1 vccd1 vccd1 _17329__1385/HI net1385 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_17_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _07498_ net335 net397 net1845 vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08837__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14510_ net1259 vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__inv_2
X_11722_ _06761_ _07153_ _07206_ net276 vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__or4b_1
XANTENNA__09880__C_N net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15490_ net1240 vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_81_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11653_ net574 _07029_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__nand2_1
X_14441_ net1272 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13043__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ net42 net41 net63 net62 vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__or4_1
XANTENNA__12397__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17160_ clknet_leaf_89_wb_clk_i _02772_ _01389_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_14372_ net1445 vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11584_ _06395_ _06397_ _06421_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13323_ net1085 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 _07749_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16111_ clknet_leaf_186_wb_clk_i _01780_ _00340_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13588__A team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10535_ _06095_ net1741 net1020 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17091_ clknet_leaf_66_wb_clk_i _02726_ _01320_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09277__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13254_ net83 team_04_WB.ADDR_START_VAL_REG\[22\] net975 vssd1 vssd1 vccd1 vccd1
+ _01652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16042_ clknet_leaf_109_wb_clk_i _01711_ _00271_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ _06036_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__nor2_1
XANTENNA__08181__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ net251 net647 vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__and2_1
X_13185_ _07621_ net379 net293 net1730 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10397_ _05728_ _05741_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08773__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12136_ net247 net2256 net511 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16944_ clknet_leaf_192_wb_clk_i _02613_ _01173_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\]
+ sky130_fd_sc_hd__dfrtp_1
X_12067_ net1949 net352 _07488_ net441 vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12857__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_53_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11018_ team_04_WB.MEM_SIZE_REG_REG\[13\] _06506_ vssd1 vssd1 vccd1 vccd1 _06507_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_159_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16875_ clknet_leaf_23_wb_clk_i _02544_ _01104_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10332__B2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15826_ clknet_leaf_92_wb_clk_i _01503_ _00053_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12609__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_142_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13282__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15757_ net1283 vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12969_ net603 _07328_ net471 net315 net1622 vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a32o_1
XANTENNA__13262__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__B net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15043__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14708_ net1225 vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__inv_2
XANTENNA__11832__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15688_ net1257 vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13034__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14639_ net1143 vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14882__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09976__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08160_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16309_ clknet_leaf_36_wb_clk_i _01978_ _00538_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14093__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ _03698_ _03699_ _03700_ _03701_ net785 net806 vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__mux4_1
X_17289_ net1345 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_31_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13337__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload30 clknet_leaf_175_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload41 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload41/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload52 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload52/X sky130_fd_sc_hd__clkbuf_8
Xclkload63 clknet_leaf_44_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11348__B1 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload74 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__clkinv_4
Xclkload85 clknet_leaf_58_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload85/Y sky130_fd_sc_hd__inv_8
Xclkload96 clknet_leaf_150_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_149_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12560__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux2_1
XANTENNA__11746__A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07944_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__nand2_8
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_166_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12848__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout373_A net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09614_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__mux2_1
XANTENNA__09650__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13273__A0 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1282_A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_174_Right_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11284__C1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09476_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08427_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__mux2_1
XANTENNA__13025__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout805_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08358_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__mux2_1
Xclkload2 clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_117_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08289_ net722 _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__or2_1
XANTENNA__10825__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10320_ _05585_ _05586_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nand2b_1
XANTENNA__09097__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net620 _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08581__A1_N net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net622 _05790_ net278 vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1206 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_2
Xfanout1215 net1220 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__buf_4
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
XANTENNA__10560__A team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1237 net1243 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_4
XANTENNA__12839__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14990_ net1197 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__inv_2
Xfanout1248 net1252 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__buf_4
Xfanout1259 net1261 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout261 _07402_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_2
Xfanout272 _07216_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13941_ _03068_ _03082_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__or2_1
Xfanout283 _05523_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_2
Xfanout294 _07683_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10314__B2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__B1 _06824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16660_ clknet_leaf_3_wb_clk_i _02329_ _00889_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\]
+ sky130_fd_sc_hd__dfrtp_1
X_13872_ net1664 net1068 _03255_ _03256_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15611_ net1114 vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__inv_2
XANTENNA__13264__A0 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _07663_ net701 net650 vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__or3b_4
X_16591_ clknet_leaf_188_wb_clk_i _02260_ _00820_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11391__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_141_Right_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15542_ net1223 vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__inv_2
X_12754_ _07479_ net344 net402 net2200 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__a22o_1
XANTENNA__08029__X _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10719__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11705_ _06271_ _06944_ _07190_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__o21ai_1
X_15473_ net1274 vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__inv_2
XANTENNA__13016__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12685_ _07445_ net2314 net478 vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__mux2_1
XANTENNA__11290__A2 _06776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_144_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17212_ net1418 _02822_ _01451_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_input91_X net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14424_ net1291 vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11636_ _05142_ net365 net361 _05141_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08904__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08669__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11578__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17143_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[8\]
+ _01372_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_14355_ net1258 vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _05446_ net467 _05470_ _05519_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__or4b_1
XFILLER_0_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13306_ net1083 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 _07732_
+ sky130_fd_sc_hd__nor2_1
X_10518_ team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] net1095 net1052 vssd1 vssd1 vccd1
+ vccd1 _06084_ sky130_fd_sc_hd__and3_1
X_14286_ _03457_ net818 _03456_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__and3b_1
X_17074_ clknet_leaf_46_wb_clk_i _00022_ _01303_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold709 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\] vssd1 vssd1
+ vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08205__A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11498_ net564 _06985_ _06986_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__a21o_1
XANTENNA__09618__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ net95 team_04_WB.MEM_SIZE_REG_REG\[4\] net984 vssd1 vssd1 vccd1 vccd1 _01666_
+ sky130_fd_sc_hd__mux2_1
X_16025_ clknet_leaf_76_wb_clk_i _00001_ _00254_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10449_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__or2_2
XFILLER_0_150_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08746__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ _07604_ net374 net291 net1619 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a22o_1
X_12119_ net2266 net354 _07514_ net455 vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11566__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ _07531_ net371 net298 net1643 vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_144_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16927_ clknet_leaf_159_wb_clk_i _02596_ _01156_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09171__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_79_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16858_ clknet_leaf_39_wb_clk_i _02527_ _01087_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_140_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16789_ clknet_leaf_33_wb_clk_i _02458_ _01018_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\]
+ sky130_fd_sc_hd__dfrtp_1
X_09330_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__mux2_1
XANTENNA__11805__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__mux2_1
XANTENNA__13007__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08212_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\]
+ net944 vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09192_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08143_ _03721_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07938__B net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08074_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__mux2_1
Xclkload130 clknet_leaf_125_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__12781__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload141 clknet_leaf_65_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload141/Y sky130_fd_sc_hd__clkinv_8
Xclkload152 clknet_leaf_92_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload152/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17328__1384 vssd1 vssd1 vccd1 vccd1 _17328__1384/HI net1384 sky130_fd_sc_hd__conb_1
Xclkload163 clknet_leaf_121_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload163/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_168_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload174 clknet_leaf_87_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload174/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_140_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09934__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_885 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09645__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11336__A3 _06824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout490_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout588_A _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10380__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\] vssd1 vssd1
+ vccd1 vccd1 net1451 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_1
Xhold25 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[19\]
+ vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 net105 vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _03535_ _03536_ _01694_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a21o_1
Xhold69 net168 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13494__B1 team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_85_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13246__A0 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout922_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08348__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ net661 _05137_ _05138_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__o21ai_2
XANTENNA__12100__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09459_ _05066_ _05067_ _05068_ _05069_ net833 net737 vssd1 vssd1 vccd1 vccd1 _05070_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12470_ net519 net601 _07471_ net428 net1731 vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__a32o_1
XANTENNA__08724__S net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13013__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11421_ net635 net634 _04724_ net632 net540 net546 vssd1 vssd1 vccd1 vccd1 _06910_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14140_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03362_
+ _03356_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.h_out sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08520__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ _06820_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__xor2_2
XFILLER_0_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12772__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _05697_ _05699_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14071_ net1490 _06088_ net1034 vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__mux2_1
XANTENNA__11938__X _07403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11283_ net568 _06694_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ net2313 net313 net383 _07481_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a22o_1
XANTENNA_input51_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _05539_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_1
XANTENNA__15854__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1001 _07685_ vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13077__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1012 net1014 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
X_10165_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] _03646_ vssd1
+ vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__xnor2_1
Xfanout1023 _06073_ vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__buf_2
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_50_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1045 net1046 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__buf_2
Xfanout1056 net1058 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_4
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13485__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _03498_ _04671_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__nand2_1
X_14973_ net1155 vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__inv_2
Xfanout1078 _03524_ vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_2
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1089 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__clkbuf_4
X_16712_ clknet_leaf_114_wb_clk_i _02381_ _00941_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\]
+ sky130_fd_sc_hd__dfrtp_1
X_13924_ _03140_ _03292_ _03132_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09290__S net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13237__A0 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16643_ clknet_leaf_125_wb_clk_i _02312_ _00872_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\]
+ sky130_fd_sc_hd__dfrtp_1
X_13855_ _03242_ _03245_ net1755 net1066 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_159_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _07349_ net2282 net322 vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__mux2_1
X_16574_ clknet_leaf_142_wb_clk_i _02243_ _00803_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\]
+ sky130_fd_sc_hd__dfrtp_1
X_13786_ net990 _03176_ _03173_ net994 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_48_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10998_ _06482_ _06486_ _06484_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15525_ net1108 vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12737_ _07462_ net336 net401 net1811 vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XANTENNA__12460__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15456_ net1212 vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11688__A_N net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12668_ net244 net2546 net477 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13004__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14407_ net1274 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12156__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _06209_ _06211_ net541 vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12212__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15387_ net1136 vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12599_ _07568_ net480 net412 net2198 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17126_ clknet_leaf_76_wb_clk_i net1556 _01355_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12763__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14338_ net1190 vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold506 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\] vssd1 vssd1
+ vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\] vssd1 vssd1
+ vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\] vssd1 vssd1
+ vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17057_ clknet_leaf_48_wb_clk_i _00035_ _01286_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold539 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\] vssd1 vssd1
+ vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
X_14269_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ _03443_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ clknet_leaf_51_wb_clk_i _01684_ _00237_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12515__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_111_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10912__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__D1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09392__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ net811 net702 _03644_ _03640_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__a22o_2
Xhold1206 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] vssd1 vssd1
+ vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__mux2_1
Xhold1228 team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\] vssd1 vssd1 vccd1
+ vccd1 net2665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08692_ _04142_ _04194_ _04249_ _04302_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and4b_1
XANTENNA__08809__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13228__A0 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_169_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09313_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12451__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09244_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08544__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09867__C _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ _03628_ _03644_ _04780_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout503_A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1245_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\]
+ net852 vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__mux2_1
XANTENNA__13951__A1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12754__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net973 _03666_ vssd1 vssd1 vccd1
+ vccd1 _03668_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_109_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09375__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12506__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__B net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout872_A net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ net726 _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _07398_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_169_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13219__A0 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _05404_ _06408_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__and3_1
XFILLER_0_86_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout925_X net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_857 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13640_ _03023_ _03029_ _03030_ team_04_WB.ADDR_START_VAL_REG\[5\] vssd1 vssd1 vccd1
+ vccd1 _03031_ sky130_fd_sc_hd__a31o_1
X_10852_ _04193_ _06301_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13571_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _05911_ net1100
+ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__mux2_1
X_10783_ net583 _06207_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__or2_4
XFILLER_0_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15310_ net1198 vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__inv_2
XANTENNA__12993__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12522_ net2302 net211 net420 vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16290_ clknet_leaf_145_wb_clk_i _01959_ _00519_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input99_A wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08307__X _03918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15849__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ net1135 vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__inv_2
X_12453_ net2527 net428 _07646_ net519 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12745__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ net540 _06869_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__or2_1
X_12384_ net261 net2616 net497 vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__mux2_1
X_15172_ net1188 vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__inv_2
XANTENNA__09610__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11953__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ team_04_WB.MEM_SIZE_REG_REG\[22\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[22\]
+ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__a22o_1
X_11335_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11828__B net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ _06279_ _06751_ _06753_ _06754_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__a211o_1
X_14054_ net33 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1
+ vccd1 vccd1 _01532_ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10217_ net620 _05821_ _05820_ net280 vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__a211o_1
X_13005_ net605 _07465_ net470 net310 net1852 vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a32o_1
XANTENNA__13170__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09141__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _06515_ _06685_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and2_1
XANTENNA__12005__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07924__A2 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _05693_ _05757_ _05694_ _05692_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o211a_1
X_10079_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__inv_2
X_14956_ net1121 vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08629__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _02958_ _02965_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__or3_1
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14887_ net1134 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_619 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327__1383 vssd1 vssd1 vccd1 vccd1 _17327__1383/HI net1383 sky130_fd_sc_hd__conb_1
X_16626_ clknet_leaf_10_wb_clk_i _02295_ _00855_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08980__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ _02863_ _03227_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16557_ clknet_leaf_29_wb_clk_i _02226_ _00786_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13769_ _06758_ net273 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__nor2_1
XANTENNA__12433__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15508_ net1235 vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12984__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ clknet_leaf_113_wb_clk_i _02157_ _00717_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12394__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15439_ net1195 vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09288__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09984__A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__A3 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__B2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold303 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\] vssd1 vssd1
+ vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_105_wb_clk_i _02744_ _01338_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[16\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold314 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\] vssd1 vssd1
+ vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\] vssd1 vssd1
+ vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold336 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\] vssd1 vssd1
+ vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\] vssd1 vssd1
+ vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09195__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold358 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\] vssd1 vssd1
+ vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\]
+ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__and3_2
XFILLER_0_110_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold369 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\] vssd1 vssd1
+ vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_863 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout805 net808 vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
XFILLER_0_68_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout816 net817 vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
XANTENNA__13161__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09862_ _04532_ _05438_ _05449_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__and4b_4
Xfanout827 net828 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11172__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout838 _03663_ vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__clkbuf_4
Xfanout849 net853 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__clkbuf_4
Xhold1003 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\] vssd1 vssd1
+ vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
X_08813_ _04420_ _04421_ _04422_ _04423_ net798 net817 vssd1 vssd1 vccd1 vccd1 _04424_
+ sky130_fd_sc_hd__mux4_1
Xhold1014 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\] vssd1 vssd1
+ vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _05386_ _05392_ _05403_ net768 vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__a22o_4
Xhold1025 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\] vssd1 vssd1
+ vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1036 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\] vssd1 vssd1
+ vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\] vssd1 vssd1
+ vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _04337_ _04343_ _04354_ net717 vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__a22o_2
Xhold1058 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\] vssd1 vssd1
+ vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08539__S net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1069 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\] vssd1 vssd1
+ vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08675_ _04282_ _04283_ _04284_ _04285_ net823 net733 vssd1 vssd1 vccd1 vccd1 _04286_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout453_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1195_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_159_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12424__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14129__X net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout718_A net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09227_ net766 _04837_ _04826_ _04820_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13968__X _03318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09279__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12727__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08109_ _03714_ _03719_ net774 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12524__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11120_ net557 net356 _06536_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold870 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\] vssd1 vssd1
+ vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold881 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\] vssd1 vssd1
+ vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _03721_ _03753_ net357 _06539_ net463 vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__o311a_1
XANTENNA__13152__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold892 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\] vssd1 vssd1
+ vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12360__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _05336_ _05341_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__nor2_1
X_14810_ net1146 vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__inv_2
XANTENNA__15136__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_A DAT_I[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ net1200 vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__inv_2
X_11953_ net1920 net528 net454 _07415_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13860__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10674__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10904_ net583 _06269_ net657 vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__o21a_1
XFILLER_0_169_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14672_ net1175 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__inv_2
X_11884_ net655 net258 vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_84_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16411_ clknet_leaf_102_wb_clk_i _02080_ _00640_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\]
+ sky130_fd_sc_hd__dfrtp_1
X_13623_ net999 _03012_ _03013_ _03007_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10835_ _06321_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__and2_1
XANTENNA__12415__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12966__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16342_ clknet_leaf_10_wb_clk_i _02011_ _00571_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\]
+ sky130_fd_sc_hd__dfrtp_1
X_13554_ _02908_ _02919_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__nor2_1
XANTENNA__11623__C1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10766_ net646 _06252_ net360 vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_41_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12505_ _07502_ net492 net427 net1693 vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a22o_1
X_16273_ clknet_leaf_171_wb_clk_i _01942_ _00502_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\]
+ sky130_fd_sc_hd__dfrtp_1
X_13485_ net706 _06651_ net273 _07697_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__o31ai_2
X_10697_ net756 _03630_ _03636_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__and3_2
XFILLER_0_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15224_ net1205 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__inv_2
XANTENNA__12718__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13915__B2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ net654 net609 net228 vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10729__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_130_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ net1233 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__inv_2
X_12367_ net241 net2599 net495 vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14106_ team_04_WB.MEM_SIZE_REG_REG\[5\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[5\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__o221a_1
XFILLER_0_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ net553 _06806_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__nor2_1
X_12298_ net2186 net501 _07593_ net450 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__a22o_1
X_15086_ net1197 vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__inv_2
XANTENNA__13679__B1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14037_ net20 net1063 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1
+ vccd1 vccd1 _01549_ sky130_fd_sc_hd__a22o_1
X_11249_ _06736_ _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13265__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15988_ clknet_leaf_79_wb_clk_i _01664_ _00217_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08359__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__B1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09044__A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14939_ net1145 vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10665__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09979__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16609_ clknet_leaf_134_wb_clk_i _02278_ _00838_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\]
+ sky130_fd_sc_hd__dfrtp_1
X_08391_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[25\] team_04_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__mux2_4
XANTENNA__14096__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10918__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12957__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09012_ net739 _04622_ net731 vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_171_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12709__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13948__B team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08822__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold100 net136 vssd1 vssd1 vccd1 vccd1 net1537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold111 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[30\] vssd1
+ vssd1 vccd1 vccd1 net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[13\] vssd1
+ vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12590__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\] vssd1 vssd1
+ vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 net113 vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08123__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\] vssd1 vssd1
+ vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[25\]
+ vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold188 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\] vssd1 vssd1
+ vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ net1056 net280 vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__nor2_4
Xfanout602 net612 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_4
Xhold199 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\] vssd1 vssd1
+ vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_2
Xfanout624 _05659_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1110_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout635 _04610_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
Xfanout646 _03589_ vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__clkbuf_4
X_09845_ _04611_ _04726_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__nand2_2
Xfanout657 _05462_ vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__buf_4
XANTENNA_input6_A DAT_I[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15952__Q team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 _07589_ vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout570_A _05251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 _07482_ vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__buf_2
XANTENNA__11484__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A _07589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09776_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12299__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout835_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10656__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__B net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10828__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08589_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13204__A team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ net58 _06156_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] net1095 net1052 vssd1 vssd1 vccd1
+ vccd1 _06106_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13270_ net97 net2644 net977 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10482_ _06051_ _06058_ _06059_ net1006 team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12221_ net228 net649 vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__and2_1
XANTENNA__10563__A team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12581__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net234 net2604 net513 vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
X_17326__1382 vssd1 vssd1 vccd1 vccd1 _17326__1382/HI net1382 sky130_fd_sc_hd__conb_1
X_11103_ net755 _06525_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_169_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_169_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16023__Q team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13125__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ clknet_leaf_139_wb_clk_i _02629_ _01189_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\]
+ sky130_fd_sc_hd__dfrtp_1
X_12083_ net2177 net352 _07496_ net437 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09563__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _06518_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__and2_1
X_15911_ clknet_leaf_123_wb_clk_i _01588_ _00138_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__dfrtp_1
X_16891_ clknet_leaf_97_wb_clk_i _02560_ _01120_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11687__A2 _06226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15862__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13085__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ clknet_leaf_90_wb_clk_i _01519_ _00069_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10895__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08179__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ net1287 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ _07637_ net472 net316 net1853 vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
XANTENNA__09501__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14724_ net1171 vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__inv_2
X_11936_ net691 _07399_ _07400_ net616 vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08907__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14655_ net1241 vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ net1941 net529 net459 _07341_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13606_ net992 _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_60_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10818_ _03975_ _04029_ _04084_ _06304_ net657 vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__o41a_1
X_14586_ net1179 vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ net704 _05810_ _07279_ _07281_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ clknet_leaf_19_wb_clk_i _01994_ _00554_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\]
+ sky130_fd_sc_hd__dfrtp_1
X_13537_ net994 _02925_ _02927_ net989 vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__o2bb2a_1
X_10749_ _06235_ _06237_ net537 vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16256_ clknet_leaf_140_wb_clk_i _01925_ _00485_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\]
+ sky130_fd_sc_hd__dfrtp_1
X_13468_ net1092 _02858_ net1044 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15207_ net1143 vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__inv_2
XANTENNA__09568__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12419_ net525 net607 _07369_ net435 net1658 vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a32o_1
X_16187_ clknet_leaf_103_wb_clk_i _01856_ _00416_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\]
+ sky130_fd_sc_hd__dfrtp_1
X_13399_ _07754_ _07824_ _07751_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__a21oi_1
Xoutput205 net205 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__11375__A1 _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12572__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15138_ net1217 vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13784__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__mux2_1
X_15069_ net1154 vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__inv_2
XANTENNA_wire257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\] vssd1 vssd1
+ vccd1 vccd1 _03506_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_155_Right_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09630_ _05237_ _05238_ _05239_ _05240_ net834 net738 vssd1 vssd1 vccd1 vccd1 _05241_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08089__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09561_ _05168_ _05169_ _05170_ _05171_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05172_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12687__X _07664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13723__S net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15504__A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__mux2_1
XANTENNA__08926__S0 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09492_ _05099_ _05100_ _05101_ _05102_ net791 net815 vssd1 vssd1 vccd1 vccd1 _05103_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08817__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08443_ _04048_ _04053_ net771 vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_A net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_173_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\]
+ net914 vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1158_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10169__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout785_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13107__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12802__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 _07661_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09383__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _07658_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
Xfanout432 _07625_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__clkbuf_8
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
Xfanout454 net457 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__clkbuf_2
X_15808__27 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__inv_2
XANTENNA_fanout952_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _06203_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__clkbuf_4
Xfanout476 _07662_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09828_ _04532_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__nand2b_2
Xfanout487 net488 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
Xfanout498 _07624_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_4
X_09759_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\]
+ net901 vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ _07497_ net336 net397 net1794 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17242__1303 vssd1 vssd1 vccd1 vccd1 _17242__1303/HI net1303 sky130_fd_sc_hd__conb_1
XFILLER_0_167_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07910__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11721_ _07140_ _07207_ _07208_ _07209_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_81_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12476__C net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14440_ net1276 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11652_ _06367_ _06865_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xor2_1
XFILLER_0_37_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11054__A0 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ net38 net37 net40 net39 vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__or4_2
XANTENNA__16018__Q net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09342__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ net1452 vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11583_ _06852_ _06949_ _07069_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__o211a_1
X_16110_ clknet_leaf_28_wb_clk_i _01779_ _00339_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08196__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13322_ net1085 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 _07748_
+ sky130_fd_sc_hd__and2_1
XANTENNA_input81_A wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09558__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17090_ clknet_leaf_75_wb_clk_i _02725_ _01319_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10534_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[22\]
+ _06094_ net1047 vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15857__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08470__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11389__A net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16041_ clknet_leaf_121_wb_clk_i _01710_ _00270_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ _06037_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__nand2_1
X_13253_ net84 team_04_WB.ADDR_START_VAL_REG\[23\] net976 vssd1 vssd1 vccd1 vccd1
+ _01653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12204_ net1977 net507 _07543_ net442 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a22o_1
X_10396_ _05618_ net617 _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__or3b_1
X_13184_ _07620_ net379 net292 net1747 vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__X _07165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ net239 net2401 net511 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XANTENNA__09293__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16943_ clknet_leaf_189_wb_clk_i _02612_ _01172_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\]
+ sky130_fd_sc_hd__dfrtp_1
X_12066_ net219 net676 vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_53_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11017_ team_04_WB.MEM_SIZE_REG_REG\[12\] _06505_ vssd1 vssd1 vccd1 vccd1 _06506_
+ sky130_fd_sc_hd__nand2b_1
X_16874_ clknet_leaf_163_wb_clk_i _02543_ _01103_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12013__A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15825_ clknet_leaf_95_wb_clk_i _01502_ _00052_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15756_ net1277 vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__inv_2
XANTENNA__12085__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ net600 _07321_ net468 net314 net1579 vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_66_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14707_ net1226 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11919_ net2175 net526 net439 _07386_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11832__A2 _07310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15687_ net1257 vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__inv_2
X_12899_ _07601_ net331 net384 net1735 vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13034__A1 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14638_ net1197 vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14569_ net1263 vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12793__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16308_ clknet_leaf_8_wb_clk_i _01977_ _00537_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08090_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\]
+ net918 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17288_ net1344 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__08225__X _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload20 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16239_ clknet_leaf_3_wb_clk_i _01908_ _00468_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload31 clknet_leaf_176_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload31/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload42 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload42/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload53 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__inv_6
Xclkload64 clknet_leaf_45_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload75 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload75/X sky130_fd_sc_hd__clkbuf_8
Xclkload86 clknet_leaf_59_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload97 clknet_leaf_151_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__11899__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11586__X _07075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10020__B2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ _04599_ _04600_ _04601_ _04602_ net797 net816 vssd1 vssd1 vccd1 vccd1 _04603_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_166_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07943_ _03552_ _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09713__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09544_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__mux2_1
XANTENNA__08547__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ net626 _05084_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__xnor2_1
X_17325__1381 vssd1 vssd1 vccd1 vccd1 _17325__1381/HI net1381 sky130_fd_sc_hd__conb_1
XANTENNA_fanout533_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1275_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08426_ net770 _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13025__A1 _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11036__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08357_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\]
+ net864 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout321_X net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__12784__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08282__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08288_ _03895_ _03896_ _03897_ _03898_ net828 net743 vssd1 vssd1 vccd1 vccd1 _03899_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _05849_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12000__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _05773_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12532__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1206 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__buf_4
Xfanout1216 net1220 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_2
Xfanout1227 net1253 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__buf_4
XANTENNA__10560__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1238 net1243 vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_4
Xfanout240 _07301_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_1
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_2
Xfanout1249 net1252 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout262 net263 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_4
X_13940_ _03085_ net1041 _03302_ net1072 net1882 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__a32o_1
Xfanout273 _07215_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout295 _07683_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11511__B2 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ _03211_ _03219_ _03254_ net1039 vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15610_ net1151 vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__inv_2
X_12822_ _07445_ net2227 net325 vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
XANTENNA__12067__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16590_ clknet_leaf_26_wb_clk_i _02259_ _00819_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15541_ net1215 vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12753_ _07478_ net345 net402 net2163 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__a22o_1
X_11704_ _07191_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15472_ net1164 vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12684_ net228 net2617 net477 vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__mux2_1
X_17211_ net1417 _02821_ _01449_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_14423_ net1291 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ net577 _06963_ _07122_ _07123_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_86_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__A1 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17142_ clknet_leaf_81_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[7\]
+ _01371_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12775__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ net1258 vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11566_ net287 _07053_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_184_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_184_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13305_ net1084 team_04_WB.MEM_SIZE_REG_REG\[25\] vssd1 vssd1 vccd1 vccd1 _07731_
+ sky130_fd_sc_hd__and2_1
X_17073_ clknet_leaf_46_wb_clk_i _00021_ _01302_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10517_ _06083_ net1507 net1022 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
X_14285_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ _03453_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__and3_1
XANTENNA__12790__X _07671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11497_ net534 _06894_ _06893_ net555 vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__o211a_1
XANTENNA__09618__S1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16024_ clknet_leaf_90_wb_clk_i _00000_ _00253_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_13236_ net96 team_04_WB.MEM_SIZE_REG_REG\[5\] net984 vssd1 vssd1 vccd1 vccd1 _01667_
+ sky130_fd_sc_hd__mux2_1
X_10448_ _06018_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_55_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_94_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11847__A team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08746__A2 _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _07603_ net368 net290 net1887 vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__a22o_1
X_10379_ _05600_ _05601_ _05619_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12118_ net221 net678 vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13098_ _07530_ net369 net298 net1837 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_144_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16926_ clknet_leaf_115_wb_clk_i _02595_ _01155_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\]
+ sky130_fd_sc_hd__dfrtp_1
X_12049_ net230 net683 vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09751__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15799__18 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__inv_2
X_16857_ clknet_leaf_152_wb_clk_i _02526_ _01086_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13273__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_159_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16788_ clknet_leaf_3_wb_clk_i _02457_ _01017_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08367__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15739_ net1287 vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__inv_2
XANTENNA__11805__A2 _07287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09987__A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__mux2_1
XANTENNA__13007__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08211_ net780 _03821_ net763 vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__o21a_1
X_09191_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12766__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08142_ _03728_ _03752_ net662 vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__mux2_2
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10645__B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08073_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
Xclkload120 clknet_leaf_138_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload120/Y sky130_fd_sc_hd__inv_6
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload131 clknet_leaf_126_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload131/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_116_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload142 clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload142/Y sky130_fd_sc_hd__inv_6
XANTENNA__12518__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload153 clknet_leaf_95_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload153/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__10792__A2 _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload164 clknet_leaf_122_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload164/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload175 clknet_leaf_88_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload175/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13956__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241__1302 vssd1 vssd1 vccd1 vccd1 _17241__1302/HI net1302 sky130_fd_sc_hd__conb_1
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09934__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1023_A _06073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _04557_ _04584_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout483_A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\] vssd1 vssd1
+ vccd1 vccd1 net1452 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 net173 vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\] vssd1 vssd1
+ vccd1 vccd1 net1474 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _03535_ _03536_ _01694_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__a21oi_1
Xhold48 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[13\]
+ vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09661__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__Y _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_X net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout748_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10600__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ net666 _03643_ _05112_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__or3_2
XFILLER_0_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08348__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout915_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09458_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1064 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08409_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\]
+ net944 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__mux2_1
XANTENNA__12527__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14308__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _06206_ _06907_ _06908_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ net706 _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__or2_1
XANTENNA__08520__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ net2650 net1056 _05897_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a21o_1
X_14070_ net1503 _06086_ net1035 vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08740__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11282_ net581 _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13182__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ net2516 net312 net380 _07480_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a22o_1
X_10233_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _05538_ vssd1
+ vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input44_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1002 _07685_ vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__buf_2
X_10164_ _05663_ _05774_ _05662_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a21o_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__clkbuf_2
Xfanout1024 _03546_ vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14131__C1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1035 _03354_ vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1046 _06177_ vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_2
X_10095_ _03498_ _04671_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nor2_1
Xfanout1057 net1058 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14972_ net1130 vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__inv_2
Xfanout1068 _07700_ vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_2
XANTENNA__13485__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 _03523_ vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09571__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__A0 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13923_ _03098_ _03141_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__and2b_1
X_16711_ clknet_leaf_168_wb_clk_i _02380_ _00940_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15870__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16642_ clknet_leaf_146_wb_clk_i _02311_ _00871_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\]
+ sky130_fd_sc_hd__dfrtp_1
X_13854_ _02853_ _03231_ _03241_ _03243_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_98_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08187__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _07340_ net2469 net325 vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
X_16573_ clknet_leaf_132_wb_clk_i _02242_ _00802_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05888_ net1100
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10997_ _06338_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__nor2_1
XANTENNA__11799__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15524_ net1183 vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12996__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12736_ _07461_ net326 net400 net2229 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XANTENNA__12460__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15455_ net1249 vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ net245 net2577 net476 vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12748__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ net1274 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_137_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11618_ _06770_ _06886_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__and2_1
XFILLER_0_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12212__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ net1142 vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ _07567_ net479 net412 net2232 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17125_ clknet_leaf_76_wb_clk_i _02760_ _01354_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_14337_ net1190 vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11549_ _07027_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\] vssd1 vssd1
+ vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09746__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold518 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\] vssd1 vssd1
+ vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ clknet_leaf_47_wb_clk_i _00034_ _01285_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold529 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\] vssd1 vssd1
+ vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14268_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ _03442_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\] vssd1 vssd1
+ vccd1 vccd1 _03446_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13268__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ clknet_leaf_50_wb_clk_i _01683_ _00236_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_150_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13173__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13219_ net83 team_04_WB.MEM_SIZE_REG_REG\[22\] net983 vssd1 vssd1 vccd1 vccd1 _01684_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11577__A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ _03361_ _03404_ _03405_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[1\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_111_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324__1380 vssd1 vssd1 vccd1 vccd1 _17324__1380/HI net1380 sky130_fd_sc_hd__conb_1
XANTENNA__12920__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10912__C _06226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1207 team_04_WB.ADDR_START_VAL_REG\[6\] vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14122__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08760_ net778 _04370_ _04365_ net762 vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__o211a_1
Xhold1218 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] vssd1 vssd1
+ vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12279__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold1229 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] vssd1
+ vssd1 vccd1 vccd1 net2666 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09481__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16909_ clknet_leaf_28_wb_clk_i _02578_ _01138_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\]
+ sky130_fd_sc_hd__dfrtp_1
X_08691_ _04273_ _04300_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_10_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13228__A1 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09312_ net629 _04919_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12987__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout329_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _03612_ _03637_ _04782_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08125_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\]
+ net852 vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__mux2_1
XANTENNA__13951__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11962__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1238_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07965__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09656__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net973 _03666_ vssd1 vssd1 vccd1
+ vccd1 _03667_ sky130_fd_sc_hd__o21a_1
XANTENNA__08560__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13164__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08266__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12911__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _04565_ _04566_ _04567_ _04568_ net837 net748 vssd1 vssd1 vccd1 vccd1 _04569_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12810__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09391__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ team_04_WB.instance_to_wrap.BUSY_O team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1
+ vccd1 _03523_ sky130_fd_sc_hd__and2b_1
XANTENNA__11934__B _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_X net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08889_ _04494_ _04499_ net772 vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__mux2_1
XANTENNA__14310__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ net552 net657 net541 vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10851_ net593 _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout918_X net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11950__A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12978__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13570_ net1093 _02960_ net1044 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10782_ net583 _06207_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__nor2_4
XFILLER_0_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_506 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09420__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ _06198_ _07657_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__nor2_8
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10566__A team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15240_ net1118 vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12452_ net600 net242 net680 vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_43_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16026__Q team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _06891_ _06888_ _06890_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__or3b_1
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15171_ net1170 vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13942__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ net250 net2433 net498 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14122_ team_04_WB.MEM_SIZE_REG_REG\[21\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[21\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__o221a_1
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11334_ net567 _06822_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__or2_1
XANTENNA__15865__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13088__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ net3 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1
+ vccd1 vccd1 _01533_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11265_ _04414_ net363 vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__nor2_1
XANTENNA__12902__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ net610 _07464_ net474 net313 net2193 vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__a32o_1
X_10216_ _05649_ _05819_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__xnor2_1
XANTENNA_input47_X net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ team_04_WB.MEM_SIZE_REG_REG\[25\] _06514_ vssd1 vssd1 vccd1 vccd1 _06685_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__12005__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10147_ _05693_ _05757_ _05694_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__o21a_1
XANTENNA__13458__A1 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14955_ net1161 vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__inv_2
X_10078_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] _04331_ vssd1
+ vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_89_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13906_ _02980_ _03280_ _02969_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a21oi_1
X_14886_ net1105 vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__inv_2
XANTENNA__12021__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13837_ _02864_ _02873_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a21oi_1
X_16625_ clknet_leaf_175_wb_clk_i _02294_ _00854_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08980__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13572__A1_N net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15332__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12969__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17240__1301 vssd1 vssd1 vccd1 vccd1 _17240__1301/HI net1301 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_139_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16556_ clknet_leaf_110_wb_clk_i _02225_ _00785_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\]
+ sky130_fd_sc_hd__dfrtp_1
X_13768_ _03157_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12433__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15507_ net1234 vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__inv_2
X_12719_ net2378 net406 net341 _07421_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16487_ clknet_leaf_165_wb_clk_i _02156_ _00716_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\]
+ sky130_fd_sc_hd__dfrtp_1
X_13699_ _03031_ _03043_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_135_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12394__C net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15438_ net1203 vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13933__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ net1137 vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11944__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold304 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[22\]
+ vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
X_17108_ clknet_leaf_64_wb_clk_i _02743_ _01337_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold315 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\] vssd1 vssd1
+ vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[1\] vssd1 vssd1
+ vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold337 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\] vssd1 vssd1
+ vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold348 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\] vssd1 vssd1
+ vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09930_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\] _05540_ vssd1
+ vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__and2_1
X_17039_ clknet_leaf_189_wb_clk_i _02708_ _01268_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10415__S net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold359 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\] vssd1 vssd1
+ vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout806 net808 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__buf_4
X_09861_ net466 _05469_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__nor2_1
Xfanout817 _03550_ vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout828 net829 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__clkbuf_8
Xfanout839 net840 vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__clkbuf_4
X_08812_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__mux2_1
X_09792_ _05397_ _05402_ net775 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__mux2_1
Xhold1004 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\] vssd1 vssd1
+ vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\] vssd1 vssd1
+ vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13525__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1026 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\] vssd1 vssd1
+ vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14110__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ _04348_ _04353_ net729 vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
Xhold1037 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\] vssd1 vssd1
+ vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\] vssd1 vssd1
+ vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\] vssd1 vssd1
+ vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_159_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1090_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10938__X _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12424__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout613_A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12975__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _04831_ _04836_ net770 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09157_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08487__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12805__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11935__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__B2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _03715_ _03716_ _03717_ _03718_ net791 net812 vssd1 vssd1 vccd1 vccd1 _03719_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09386__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08290__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ _04668_ _04697_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout982_A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Right_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13137__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ net1079 net1028 net1024 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__a31oi_4
XANTENNA__12106__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\] vssd1 vssd1
+ vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11010__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\] vssd1 vssd1
+ vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap590 _04812_ vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold882 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\] vssd1 vssd1
+ vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _03721_ _03753_ net360 vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__a21o_1
Xhold893 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\] vssd1 vssd1
+ vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13636__S net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08022__C net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _05404_ _05408_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__nand2_1
XANTENNA__11945__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__X _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14740_ net1208 vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__inv_2
X_11952_ net654 net223 vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__and2_1
XANTENNA__13860__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _06390_ _06391_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10674__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ net1140 vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__inv_2
X_11883_ net690 _06879_ _07355_ net613 vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__o211a_2
X_16410_ clknet_leaf_38_wb_clk_i _02079_ _00639_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_84_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ net991 _03011_ _03009_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10834_ net644 _06320_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12415__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13612__B2 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09150__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16341_ clknet_leaf_37_wb_clk_i _02010_ _00570_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\]
+ sky130_fd_sc_hd__dfrtp_1
X_13553_ _02922_ _02933_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__nor3_1
XFILLER_0_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10765_ _05450_ net467 _05470_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__or3_2
XANTENNA__14991__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12504_ _07501_ net488 net427 net1661 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
X_16272_ clknet_leaf_190_wb_clk_i _01941_ _00501_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__and2b_1
X_10696_ net905 net752 vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_4
XANTENNA_output198_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15223_ net1230 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ net2255 net434 _07638_ net524 vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11926__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ net1246 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ net226 net2355 net495 vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14105_ team_04_WB.MEM_SIZE_REG_REG\[4\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__a22o_1
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13128__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11317_ net530 _06527_ _06528_ _06805_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__a31oi_1
X_15085_ net1152 vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__inv_2
X_12297_ net213 net670 vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__and2_1
XANTENNA__13679__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ net21 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1
+ vccd1 vccd1 _01550_ sky130_fd_sc_hd__o22a_1
X_11248_ _06548_ _06551_ net530 vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11179_ net566 _06666_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ clknet_leaf_72_wb_clk_i _01663_ _00216_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12103__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14938_ net1151 vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__inv_2
XANTENNA__11311__C1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09612__X _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10665__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ net1211 vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16608_ clknet_leaf_140_wb_clk_i _02277_ _00837_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08390_ net766 _04000_ _03989_ _03988_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08375__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12957__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16539_ clknet_leaf_98_wb_clk_i _02208_ _00768_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_154_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09995__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09011_ _04618_ _04619_ _04620_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o22a_1
XFILLER_0_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_171_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_171_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11917__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold101 net163 vssd1 vssd1 vccd1 vccd1 net1538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\] vssd1 vssd1
+ vccd1 vccd1 net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\] vssd1 vssd1
+ vccd1 vccd1 net1560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13119__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14316__C1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold134 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[31\] vssd1
+ vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold145 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[29\]
+ vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold156 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\] vssd1 vssd1
+ vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 net116 vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net280 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__inv_2
Xhold178 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\] vssd1 vssd1
+ vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[6\] vssd1 vssd1
+ vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13964__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout603 net604 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__buf_2
Xfanout614 _06193_ vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__buf_4
XANTENNA_fanout396_A _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 _05276_ vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12342__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout636 _04501_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12360__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _04726_ _05453_ _05454_ _05444_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__o2bb2a_1
Xfanout647 _07520_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_8
Xfanout658 _05461_ vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1103_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 _07589_ vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11484__B _06972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09235__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ net775 _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout563_A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ net723 _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12645__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08657_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout730_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout828_A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08285__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ _04195_ _04196_ _04197_ _04198_ net783 net805 vssd1 vssd1 vccd1 vccd1 _04199_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10408__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11605__B1 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17303__1359 vssd1 vssd1 vccd1 vccd1 _17303__1359/HI net1359 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_12_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15700__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11081__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _06105_ net1536 net1021 vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08017__C net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09209_ net771 _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _06006_ _06057_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12535__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ net2074 net509 _07551_ net455 vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a22o_1
XANTENNA__10563__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12151_ net261 net2472 net513 vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_783 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11102_ _05473_ _06538_ _06542_ _06590_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__or4b_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ net246 net676 vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__and2_1
Xhold690 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\] vssd1 vssd1
+ vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11033_ team_04_WB.MEM_SIZE_REG_REG\[29\] _06517_ team_04_WB.MEM_SIZE_REG_REG\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__o21ai_1
X_15910_ clknet_leaf_12_wb_clk_i _01587_ _00137_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10344__B1 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16890_ clknet_leaf_39_wb_clk_i _02559_ _01119_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12884__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ clknet_leaf_87_wb_clk_i _01518_ _00068_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_138_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_86_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15772_ net1287 vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__inv_2
X_12984_ _07636_ net473 net316 net1690 vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__a22o_1
XANTENNA__12636__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11935_ net905 _03630_ _05961_ _05959_ net756 vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__o32a_1
X_14723_ net1170 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11844__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14654_ net1217 vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08195__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11866_ net655 net244 vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13605_ _07802_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10817_ _04029_ _04084_ _06304_ net657 vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__o31a_1
X_14585_ net1186 vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ net686 _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13536_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _05854_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16324_ clknet_leaf_167_wb_clk_i _01993_ _00553_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08923__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ net592 net549 _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ clknet_leaf_156_wb_clk_i _01924_ _00484_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13467_ _07874_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10679_ net2465 net1017 net1013 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1
+ vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_531 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15206_ net1104 vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12418_ net525 net611 _07363_ net435 net1580 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a32o_1
XANTENNA__11569__B _07057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16186_ clknet_leaf_44_wb_clk_i _01855_ _00415_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\]
+ sky130_fd_sc_hd__dfrtp_1
X_13398_ _07822_ _07823_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput206 net206 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_112_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15137_ net1169 vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ net231 net670 vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08871__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09754__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15068_ net1130 vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__inv_2
XANTENNA__08528__A0 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ _05466_ _03345_ _07694_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__a21o_1
XANTENNA__12324__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07890_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\] vssd1 vssd1
+ vccd1 vccd1 _03505_ sky130_fd_sc_hd__inv_2
XANTENNA__12875__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11872__X _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__mux2_1
XANTENNA__13338__C_N team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12627__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08511_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\]
+ net846 vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__mux2_1
X_09491_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__mux2_1
XANTENNA__08926__S1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_43_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13305__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08442_ _04049_ _04050_ _04051_ _04052_ net785 net806 vssd1 vssd1 vccd1 vccd1 _04053_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10648__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13052__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11063__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10810__A1 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout311_A _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout409_A _07661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09664__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _07669_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_6
Xfanout411 _07661_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout778_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _07658_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_6
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout433 _07625_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_4
Xfanout444 _07252_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12866__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout455 net456 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_4
Xfanout466 _05465_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
Xfanout477 _07662_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_6
X_09827_ _04755_ _04978_ _05195_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__and4_1
Xfanout488 net491 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_4
XANTENNA_fanout945_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 net500 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__clkbuf_8
X_09758_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12618__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _04316_ _04317_ _04318_ _04319_ net787 net810 vssd1 vssd1 vccd1 vccd1 _04320_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_61_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _05296_ _05297_ _05298_ _05299_ net834 net746 vssd1 vssd1 vccd1 vccd1 _05300_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10839__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08309__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11651_ _07136_ _07138_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout900_X net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13043__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ net101 net68 net102 vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11054__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14370_ net1468 vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08743__S net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09342__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ _06847_ _06886_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ net1085 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 _07747_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06094_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16040_ clknet_leaf_110_wb_clk_i _01709_ _00269_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_13252_ net85 team_04_WB.ADDR_START_VAL_REG\[24\] net975 vssd1 vssd1 vccd1 vccd1
+ _01654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10464_ _06041_ _06042_ _06039_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__a21o_1
XANTENNA_input74_A wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12203_ net253 net647 vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ _07619_ net376 net292 net2029 vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a22o_1
X_10395_ _05605_ _05606_ _05617_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__or3_1
XANTENNA__09574__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ net241 net2477 net511 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15873__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10513__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16942_ clknet_leaf_42_wb_clk_i _02611_ _01171_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\]
+ sky130_fd_sc_hd__dfrtp_1
X_12065_ net2023 net354 _07487_ net450 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
XANTENNA__08605__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ team_04_WB.MEM_SIZE_REG_REG\[10\] _06504_ team_04_WB.MEM_SIZE_REG_REG\[11\]
+ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__a21oi_2
X_16873_ clknet_leaf_123_wb_clk_i _02542_ _01102_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14059__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12013__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15824_ clknet_leaf_97_wb_clk_i _01501_ _00051_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_149_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12609__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08908__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15755_ net1275 vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__inv_2
X_12967_ _07633_ net468 net314 net1820 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ net651 net253 vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__and2_1
X_14706_ net1237 vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__inv_2
XANTENNA__12490__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15686_ net1256 vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__inv_2
X_12898_ _07600_ net328 net384 net1739 vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ net689 _06729_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__or2_1
X_14637_ net1210 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__inv_2
XFILLER_0_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13034__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14568_ net1264 vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__inv_2
XANTENNA__08653__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_109_Left_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16307_ clknet_leaf_182_wb_clk_i _01976_ _00536_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13519_ _02908_ _02909_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14499_ net1263 vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__inv_2
X_17287_ net1343 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_141_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload10 clknet_leaf_182_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_152_160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload21 clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/X sky130_fd_sc_hd__clkbuf_8
Xclkload32 clknet_leaf_177_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload32/X sky130_fd_sc_hd__clkbuf_8
X_16238_ clknet_leaf_31_wb_clk_i _01907_ _00467_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[211\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload43 clknet_leaf_164_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__12545__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload54 clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__inv_6
XANTENNA__11348__A2 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13742__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload65 clknet_leaf_46_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_77_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload76 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload76/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload87 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ clknet_leaf_120_wb_clk_i _01838_ _00398_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_152_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload98/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09484__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_188_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08991_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07942_ team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] net1078 net1030 net1026 vssd1
+ vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__or4_4
XANTENNA__10308__B1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12848__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17302__1358 vssd1 vssd1 vccd1 vccd1 _17302__1358/HI net1358 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_3_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4__f_wb_clk_i_X clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09612_ net731 _03722_ net700 _03637_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a22o_2
XTAP_TAPCELL_ROW_3_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09543_ net775 _05147_ _05153_ net763 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__o211a_1
XANTENNA__11808__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09474_ net626 _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__and2_1
X_08425_ _04032_ _04033_ _04034_ _04035_ net785 net806 vssd1 vssd1 vccd1 vccd1 _04036_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_148_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13025__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A _06195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1268_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09659__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08356_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11789__A1_N net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload4 clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__inv_6
XFILLER_0_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08287_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout314_X net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13201__C net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout895_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12536__A1 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12813__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10180_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13992__X _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1254 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__buf_2
X_15787__6 clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__inv_2
Xfanout1217 net1219 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_4
Xfanout1228 net1230 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
XANTENNA__12114__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _07426_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12839__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout241 _07295_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_2
XANTENNA__10560__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1239 net1242 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout263 _07234_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
Xfanout274 net275 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__buf_6
XANTENNA__11511__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ _03219_ _03254_ _03211_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08738__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ net228 net2611 net324 vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
XANTENNA__10569__A team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15540_ net1235 vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__inv_2
X_12752_ _07477_ net351 net402 net2348 vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12472__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11703_ _03946_ _03975_ _06257_ _06279_ _06947_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__a32o_1
X_15471_ net1195 vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12683_ net222 net2603 net477 vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__mux2_1
XANTENNA__13016__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17210_ net1416 _02820_ _01447_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_14422_ net1283 vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__inv_2
XANTENNA__09569__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11634_ net555 _07002_ net569 vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15868__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17141_ clknet_leaf_81_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[6\]
+ _01370_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_14353_ net1258 vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10508__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ _06885_ _06923_ _07049_ _06278_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire642 _03945_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08045__Y _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13304_ net1082 team_04_WB.MEM_SIZE_REG_REG\[25\] vssd1 vssd1 vccd1 vccd1 _07730_
+ sky130_fd_sc_hd__nor2_1
X_17072_ clknet_leaf_46_wb_clk_i _00020_ _01301_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10516_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[28\]
+ _06082_ net1049 vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_98_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input77_X net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14284_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\]
+ _03452_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[23\] vssd1 vssd1
+ vccd1 vccd1 _03456_ sky130_fd_sc_hd__a31o_1
XANTENNA_output180_A net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11496_ net634 net632 net630 net628 net546 net539 vssd1 vssd1 vccd1 vccd1 _06985_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12527__A1 _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ net97 team_04_WB.MEM_SIZE_REG_REG\[6\] net984 vssd1 vssd1 vccd1 vccd1 _01668_
+ sky130_fd_sc_hd__mux2_1
X_16023_ clknet_leaf_77_wb_clk_i _01695_ _00252_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.BUSY_O
+ sky130_fd_sc_hd__dfrtp_4
X_10447_ _06017_ _06020_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__and2b_1
XFILLER_0_27_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08826__S0 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14504__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13166_ _07602_ net367 net290 net1744 vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__a22o_1
X_10378_ net2660 _05964_ net1076 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XANTENNA__10751__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_153_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_153_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12117_ net2594 net354 _07513_ net456 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13097_ _07529_ net367 net298 net1895 vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09156__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16925_ clknet_leaf_132_wb_clk_i _02594_ _01154_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\]
+ sky130_fd_sc_hd__dfrtp_1
X_12048_ net2337 net517 _07477_ net452 vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a22o_1
XANTENNA__09251__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08903__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16856_ clknet_leaf_148_wb_clk_i _02525_ _01085_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10710__B1 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16787_ clknet_leaf_184_wb_clk_i _02456_ _01016_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\]
+ sky130_fd_sc_hd__dfrtp_1
X_13999_ net1531 net1069 _03334_ net265 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__a22o_1
X_15738_ net1264 vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12463__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15669_ net1282 vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08210_ _03817_ _03818_ _03819_ _03820_ net791 net802 vssd1 vssd1 vccd1 vccd1 _03821_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09479__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12766__A1 _07493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ net718 _03751_ _03740_ _03734_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__o2bb2a_2
X_17339_ net1395 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11103__A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload110 clknet_leaf_159_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload110/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_70_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08072_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload121 clknet_leaf_139_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_116_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload132 clknet_leaf_127_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__clkinv_2
Xclkload143 clknet_leaf_67_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload143/Y sky130_fd_sc_hd__clkinv_8
Xclkload154 clknet_leaf_96_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload154/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_144_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10942__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload165 clknet_leaf_123_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload165/X sky130_fd_sc_hd__clkbuf_4
Xclkload176 clknet_leaf_89_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload176/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09508__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_126_Left_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08974_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1016_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\] vssd1 vssd1
+ vccd1 vccd1 net1453 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07925_ net1101 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\]
+ net1080 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__mux2_1
Xhold27 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13972__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[23\]
+ vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08558__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout643_A _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ _05119_ _05125_ _05136_ net718 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__a22o_2
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_135_Left_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout810_A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12808__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout908_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_X net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09389__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08408_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__mux2_1
XANTENNA__08293__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10217__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14308__B net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11965__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11350_ net463 _06821_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_105_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12509__A1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10301_ _05891_ _05893_ _05896_ net278 net1075 vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12543__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11281_ net576 _06691_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08808__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13020_ _06189_ _07250_ _07665_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor3_4
X_10232_ net621 _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 net1005 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__clkbuf_4
X_10163_ _05665_ _05773_ _05666_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a21bo_1
Xfanout1014 _06178_ vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_2
XANTENNA__10940__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08041__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1025 _03546_ vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14131__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1047 net1050 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__clkbuf_4
X_10094_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] _04728_ vssd1
+ vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__nand2_1
X_14971_ net1136 vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__inv_2
XANTENNA__13485__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 _03526_ vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1069 net1070 vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16710_ clknet_leaf_22_wb_clk_i _02379_ _00939_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\]
+ sky130_fd_sc_hd__dfrtp_1
X_13922_ _03288_ _03291_ net104 net1071 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11496__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12693__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16641_ clknet_leaf_134_wb_clk_i _02310_ _00870_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13853_ net1 net1072 vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12804_ net245 net2627 net323 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__mux2_1
XANTENNA__09536__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16572_ clknet_leaf_126_wb_clk_i _02241_ _00801_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\]
+ sky130_fd_sc_hd__dfrtp_1
X_13784_ net1002 _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10996_ _06334_ _06483_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__nand2_1
XANTENNA__11799__A2 _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12996__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15523_ net1182 vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ _07460_ net326 net400 net2089 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15454_ net1236 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__inv_2
X_12666_ net260 net2318 net476 vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13945__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14405_ net1274 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__inv_2
X_11617_ _05404_ net533 _06253_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__o21a_1
X_17301__1357 vssd1 vssd1 vccd1 vccd1 _17301__1357/HI net1357 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_137_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _07566_ net481 net412 net1862 vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22o_1
X_15385_ net1250 vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17124_ clknet_leaf_65_wb_clk_i _02759_ _01353_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_14336_ net1190 vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11548_ net286 _07034_ _07036_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__or3_2
XANTENNA__08931__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold508 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] vssd1 vssd1
+ vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11858__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14267_ net1915 _03443_ _03445_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__a21oi_1
X_17055_ clknet_leaf_48_wb_clk_i _00033_ _01284_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold519 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\] vssd1 vssd1
+ vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ _05464_ _06535_ _06967_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__o21a_1
X_16006_ clknet_leaf_51_wb_clk_i _01682_ _00235_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_13218_ net84 team_04_WB.MEM_SIZE_REG_REG\[23\] net983 vssd1 vssd1 vccd1 vccd1 _01685_
+ sky130_fd_sc_hd__mux2_1
X_14198_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1090
+ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07927__A1 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12920__A1 _07622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ _07583_ net378 net296 net2114 vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09129__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14122__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1208 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\] vssd1 vssd1
+ vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1219 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] vssd1 vssd1
+ vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12684__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16908_ clknet_leaf_119_wb_clk_i _02577_ _01137_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\]
+ sky130_fd_sc_hd__dfrtp_1
X_08690_ _04300_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__inv_2
X_16839_ clknet_leaf_166_wb_clk_i _02508_ _01068_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_89 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09998__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09311_ net628 _04919_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13936__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09173_ net905 _03612_ _03624_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__and3_2
XFILLER_0_56_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout224_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08124_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13951__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[23\] net1009
+ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__or2_1
XANTENNA__12363__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08266__S1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13983__A _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10922__B1 _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__A team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__15971__Q team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout760_A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ _04495_ _04496_ _04497_ _04498_ net788 net809 vssd1 vssd1 vccd1 vccd1 _04499_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13207__B _06145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15703__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _04139_ _06302_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12978__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09701__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09509_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ net584 net466 _06251_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__or3_1
XANTENNA__10847__A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12520_ net700 _07517_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__or2_2
XFILLER_0_136_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07946__A_N net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ net519 net600 _07456_ net428 net2041 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_43_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11402_ net582 _06603_ _06610_ _06886_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__a22o_1
X_15170_ net1217 vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__inv_2
XANTENNA__11402__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ net252 net2470 net496 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14121_ team_04_WB.MEM_SIZE_REG_REG\[20\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[20\]
+ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__a22o_1
XFILLER_0_50_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11953__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _06801_ _06806_ net554 vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14052_ net4 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1
+ vccd1 vccd1 _01534_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_91_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11264_ _04385_ _04413_ _06257_ _06752_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ net604 _07463_ net470 net311 net1742 vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a32o_1
XANTENNA__12902__A1 _07604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ net620 _05818_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nor2_1
XANTENNA__11965__X _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11195_ _06681_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10913__B1 _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08582__A1 _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _05696_ _05756_ _05695_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10077_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _04219_ vssd1
+ vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__xnor2_1
X_14954_ net1105 vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08334__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ _02981_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nand2_1
X_14885_ net1111 vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__inv_2
XANTENNA__12021__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16624_ clknet_leaf_190_wb_clk_i _02293_ _00853_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15613__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ team_04_WB.ADDR_START_VAL_REG\[29\] _02856_ _02862_ vssd1 vssd1 vccd1 vccd1
+ _03227_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12418__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12969__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08098__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16555_ clknet_leaf_30_wb_clk_i _02224_ _00784_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\]
+ sky130_fd_sc_hd__dfrtp_1
X_13767_ team_04_WB.ADDR_START_VAL_REG\[19\] _03156_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_139_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10979_ _06466_ _06467_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__nand2_1
XANTENNA__13091__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15506_ net1247 vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__inv_2
X_12718_ net2084 net406 net342 _07415_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ clknet_leaf_17_wb_clk_i _02155_ _00715_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\]
+ sky130_fd_sc_hd__dfrtp_1
X_13698_ team_04_WB.ADDR_START_VAL_REG\[5\] _03023_ _03029_ _03030_ vssd1 vssd1 vccd1
+ vccd1 _03089_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15437_ net1143 vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12649_ _07620_ net489 net410 net1713 vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09757__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15368_ net1125 vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12691__B net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13279__S _05525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17107_ clknet_leaf_63_wb_clk_i _02742_ _01336_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_14319_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[27\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[26\] net1091
+ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__mux2_1
Xhold305 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\] vssd1 vssd1
+ vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold316 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\] vssd1 vssd1
+ vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ net1168 vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold327 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold338 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\] vssd1 vssd1
+ vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17038_ clknet_leaf_28_wb_clk_i _02707_ _01267_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold349 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\] vssd1 vssd1
+ vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14899__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11875__X _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _05439_ _05449_ net466 _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and4_1
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout807 net808 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_2
XFILLER_0_110_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout818 net821 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08897__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10904__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__clkbuf_8
X_08811_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\]
+ net972 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__mux2_1
X_09791_ _05398_ _05399_ _05400_ _05401_ net794 net814 vssd1 vssd1 vccd1 vccd1 _05402_
+ sky130_fd_sc_hd__mux4_1
Xhold1005 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\] vssd1 vssd1
+ vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\] vssd1 vssd1
+ vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _04349_ _04350_ _04351_ _04352_ net827 net744 vssd1 vssd1 vccd1 vccd1 _04353_
+ sky130_fd_sc_hd__mux4_1
Xhold1027 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\] vssd1 vssd1
+ vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12657__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1038 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\] vssd1 vssd1
+ vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1049 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\] vssd1 vssd1
+ vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_139_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12121__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08673_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13082__A0 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09225_ _04832_ _04833_ _04834_ _04835_ net784 net805 vssd1 vssd1 vccd1 vccd1 _04836_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_20_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13978__A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1035 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout606_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17344__1400 vssd1 vssd1 vccd1 vccd1 _17344__1400/HI net1400 sky130_fd_sc_hd__conb_1
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12188__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09156_ net772 _04766_ net761 vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08571__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08487__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09087_ _04697_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net974 _03647_ vssd1 vssd1 vccd1
+ vccd1 _03649_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold850 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\] vssd1 vssd1
+ vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11148__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12106__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\] vssd1 vssd1
+ vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11785__X _07271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__B _06498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold872 team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\] vssd1 vssd1
+ vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap591 _04384_ vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__buf_4
Xhold883 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\] vssd1 vssd1
+ vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12821__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold894 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\] vssd1 vssd1
+ vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _05609_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__nand2_1
XANTENNA__08022__D net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09989_ _05598_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12648__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17300__1356 vssd1 vssd1 vccd1 vccd1 _17300__1356/HI net1356 sky130_fd_sc_hd__conb_1
XANTENNA__13845__C1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11951_ net695 _07075_ _07413_ net616 vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_118_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13647__A1_N net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11961__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _05056_ _06389_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__and2_1
X_11882_ net687 _07354_ _07352_ _07351_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a211o_1
XANTENNA__10674__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ net1197 vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13621_ _06175_ _03011_ _03010_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__a21oi_1
X_10833_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13073__A0 _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16340_ clknet_leaf_8_wb_clk_i _02009_ _00569_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11623__A1 _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13552_ _02941_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10764_ _05449_ _05464_ _05469_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and3_1
XANTENNA__08047__A team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_165_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _07500_ net484 net425 net1753 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
X_13483_ _02865_ _02869_ _02872_ team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1
+ vccd1 _02874_ sky130_fd_sc_hd__a31o_1
X_16271_ clknet_leaf_3_wb_clk_i _01940_ _00500_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ _03608_ _03630_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__nor2_2
XFILLER_0_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15222_ net1224 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__inv_2
XANTENNA__09577__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12434_ net654 net608 net221 vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__and3_1
XANTENNA__15876__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13400__B team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12365_ net227 net2317 net496 vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__mux2_1
X_15153_ net1272 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__inv_2
XANTENNA__10516__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14104_ team_04_WB.MEM_SIZE_REG_REG\[3\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[3\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__o221a_1
X_11316_ net538 _06561_ _06563_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__and3_1
X_15084_ net1119 vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__inv_2
X_12296_ net2169 net500 _07592_ net448 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a22o_1
XANTENNA__13679__A2 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14035_ net22 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1
+ vccd1 vccd1 _01551_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _06544_ _06549_ net530 vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12887__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14512__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08555__A1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ net566 _06529_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__nand2_1
X_10129_ _05733_ _05739_ _05732_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__a21o_1
XANTENNA__12639__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15986_ clknet_leaf_72_wb_clk_i _01662_ _00215_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_69_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12103__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08307__B2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ net1241 vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11871__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11862__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08656__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14868_ net1214 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__inv_2
X_16607_ clknet_leaf_156_wb_clk_i _02276_ _00836_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\]
+ sky130_fd_sc_hd__dfrtp_1
X_13819_ _03201_ _03205_ _03208_ team_04_WB.ADDR_START_VAL_REG\[25\] vssd1 vssd1 vccd1
+ vccd1 _03210_ sky130_fd_sc_hd__a31o_1
X_14799_ net1143 vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16538_ clknet_leaf_38_wb_clk_i _02207_ _00767_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12811__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16469_ clknet_leaf_35_wb_clk_i _02138_ _00698_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09010_ _03506_ net1008 net1007 _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__a311o_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08391__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_94_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11917__A2 _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold102 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[10\]
+ vssd1 vssd1 vccd1 vccd1 net1539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12207__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold113 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\] vssd1 vssd1
+ vccd1 vccd1 net1550 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\] vssd1 vssd1
+ vccd1 vccd1 net1561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 net142 vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\] vssd1 vssd1
+ vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_04_WB.instance_to_wrap.final_design.uart.working_data\[1\] vssd1 vssd1
+ vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _05471_ _05473_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__nor3_4
Xhold179 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\] vssd1 vssd1
+ vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__buf_2
Xfanout615 _06192_ vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_8
Xfanout626 _05056_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12342__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _04611_ _04669_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout648 _07520_ vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__buf_2
Xfanout659 _05461_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_A _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout389_A _07673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09774_ _05381_ _05382_ _05383_ _05384_ net794 net814 vssd1 vssd1 vccd1 vccd1 _05385_
+ sky130_fd_sc_hd__mux4_1
X_08725_ _04332_ _04333_ _04334_ _04335_ net829 net735 vssd1 vssd1 vccd1 vccd1 _04336_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13980__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11853__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
XANTENNA__08566__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__B2 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
XANTENNA__13055__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12802__A0 _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout511_X net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12816__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1253_X net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13358__A1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _04815_ _04816_ _04817_ _04818_ net784 net805 vssd1 vssd1 vccd1 vccd1 _04819_
+ sky130_fd_sc_hd__mux4_1
X_10480_ _06006_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09139_ _04746_ _04747_ _04748_ _04749_ net834 net746 vssd1 vssd1 vccd1 vccd1 _04750_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12030__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__A team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12581__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ net250 net2478 net514 vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout978_X net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _06271_ _06589_ _06567_ net585 vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__a2bb2o_1
X_12081_ net1908 net352 _07495_ net436 vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a22o_1
XANTENNA__12551__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12869__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10860__A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\] vssd1 vssd1
+ vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\] vssd1 vssd1
+ vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _06499_ _06519_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__and2_1
XANTENNA__10344__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ clknet_leaf_87_wb_clk_i _01517_ _00067_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15771_ net1287 vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _07635_ net472 net316 net1688 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a22o_1
XANTENNA__12097__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14722_ net1218 vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__inv_2
X_11934_ _07238_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_178_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_178_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13046__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14653_ net1149 vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__inv_2
X_11865_ net613 _07338_ _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13604_ _07781_ _07783_ _07801_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_107_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10816_ _04084_ net657 _06304_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a21oi_1
X_14584_ net1179 vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__inv_2
X_11796_ team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] net270 net268 vssd1 vssd1 vccd1
+ vccd1 _07280_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16323_ clknet_leaf_121_wb_clk_i _01992_ _00552_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ net1092 _02925_ net1043 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11072__A2 _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10747_ net593 net543 vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16254_ clknet_leaf_142_wb_clk_i _01923_ _00483_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\]
+ sky130_fd_sc_hd__dfrtp_1
X_13466_ _07867_ _07870_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__nor2_1
X_10678_ net1620 net1017 net1013 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1
+ vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15205_ net1109 vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08225__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net522 net610 _07357_ net433 net1736 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a32o_1
XFILLER_0_23_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16185_ clknet_leaf_175_wb_clk_i _01854_ _00414_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\]
+ sky130_fd_sc_hd__dfrtp_1
X_13397_ team_04_WB.MEM_SIZE_REG_REG\[16\] _07753_ _07754_ vssd1 vssd1 vccd1 vccd1
+ _07823_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08999__X _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12027__A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput207 net207 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XANTENNA__08776__A1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ net1211 vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__inv_2
XANTENNA__12572__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ net2105 net501 _07618_ net453 vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_178_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08871__S1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11866__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ net2463 net505 _07582_ net454 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__a22o_1
X_15067_ net1113 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__inv_2
XANTENNA__08528__A1 _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12324__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _05338_ _07235_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_147_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09770__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15969_ clknet_leaf_50_wb_clk_i _01645_ _00198_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08510_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__mux2_1
XANTENNA__15073__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09490_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08386__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08441_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13037__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08139__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_173_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_173_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10945__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12012__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout304_A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12371__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 _07669_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_4
Xfanout412 net415 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__clkbuf_8
Xfanout423 _07658_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_4
Xfanout434 _07625_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_4
XANTENNA__08150__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_A _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout445 net446 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_2
Xfanout456 net457 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
X_09826_ _05252_ _05312_ _05380_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__nor4_1
Xfanout467 _05465_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_1
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout478 _07662_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_4
Xfanout489 net491 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09680__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13276__A0 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout938_A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11826__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08708_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\]
+ net937 vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
XANTENNA__12400__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08296__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__mux2_1
XANTENNA__13028__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11650_ _07011_ _07024_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15711__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10601_ _06139_ net1618 net1022 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ net576 _06896_ _07065_ _06277_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__o211a_1
XANTENNA__10855__A _04166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12251__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12546__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ net1085 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 _07746_
+ sky130_fd_sc_hd__nor2_1
X_10532_ _06093_ net1559 net1020 vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10463_ _06033_ _06040_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__xnor2_1
X_13251_ net86 team_04_WB.ADDR_START_VAL_REG\[25\] net976 vssd1 vssd1 vccd1 vccd1
+ _01655_ sky130_fd_sc_hd__mux2_1
X_12202_ net2295 net507 _07542_ net439 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a22o_1
X_13182_ _07618_ net378 net292 net1776 vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a22o_1
XANTENNA_input67_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ net2664 _05978_ net1076 vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ net226 net2596 net511 vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10590__A team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12306__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16941_ clknet_leaf_42_wb_clk_i _02610_ _01170_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\]
+ sky130_fd_sc_hd__dfrtp_1
X_12064_ net215 net678 vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__and2_2
XANTENNA__08605__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14997__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ team_04_WB.MEM_SIZE_REG_REG\[9\] _06503_ vssd1 vssd1 vccd1 vccd1 _06504_
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_53_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16872_ clknet_leaf_116_wb_clk_i _02541_ _01101_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout990 net991 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09590__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__A0 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15823_ clknet_leaf_92_wb_clk_i _01500_ _00050_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11817__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15754_ net1275 vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _07632_ net469 net314 net1779 vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14705_ net1274 vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ net691 _06954_ _07384_ net614 vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__o211a_4
XTAP_TAPCELL_ROW_16_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__B1 net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15685_ net1256 vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12897_ _07599_ net329 net384 net1849 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14636_ net1128 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__inv_2
X_11848_ net268 _07324_ net687 vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08446__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14567_ net1185 vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11779_ net2327 net528 net450 _07265_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ clknet_leaf_9_wb_clk_i _01975_ _00535_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\]
+ sky130_fd_sc_hd__dfrtp_1
X_13518_ _02901_ _02907_ team_04_WB.ADDR_START_VAL_REG\[23\] vssd1 vssd1 vccd1 vccd1
+ _02909_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17286_ net1342 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
X_14498_ net1263 vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16237_ clknet_leaf_41_wb_clk_i _01906_ _00466_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload11 clknet_leaf_185_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinv_2
X_13449_ _07727_ _07867_ _07873_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_113_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload22 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload33 clknet_leaf_178_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__clkinv_2
Xclkbuf_leaf_75_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload44 clknet_leaf_165_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload44/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_140_334 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload55 clknet_leaf_32_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload66 clknet_leaf_47_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_6
X_16168_ clknet_leaf_110_wb_clk_i _01837_ _00397_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload77 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload77/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload88 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__inv_6
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload99 clknet_leaf_153_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload99/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_149_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ net1140 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16099_ clknet_leaf_117_wb_clk_i _01768_ _00328_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_08990_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__mux2_1
XANTENNA__09066__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ net1080 net1029 net1025 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_166_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11883__X _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\] net1010
+ _05220_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_3_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09542_ net780 _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or2_1
X_15813__32 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__inv_2
XFILLER_0_148_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ net665 _05083_ _05059_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_116_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12481__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_A _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__mux2_1
XANTENNA__08844__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08355_ _03962_ _03963_ _03964_ _03965_ net828 net743 vssd1 vssd1 vccd1 vccd1 _03966_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12366__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12233__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_A _07658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10244__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout519_A net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12784__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload5 clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__inv_6
XANTENNA__13981__A1 _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08286_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13986__A _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout790_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1207 net1209 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_4
Xfanout220 _07271_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net1219 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__buf_4
XANTENNA__12889__X _07674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1229 net1230 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__buf_2
XANTENNA__12114__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__buf_2
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 _07295_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_1
XANTENNA__15706__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout253 _07385_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_2
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14610__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout286 _06206_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_2
X_09809_ net730 _05419_ net714 vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__o21a_1
Xfanout297 _07683_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_4
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ net221 net2455 net325 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08676__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12751_ _07476_ net342 net402 net2072 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__a22o_1
XANTENNA__12472__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11702_ _03977_ net363 net362 _03976_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08771__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15470_ net1203 vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12682_ net229 net2571 net477 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__mux2_1
XANTENNA__08607__X _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14421_ net1283 vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11633_ net532 _07046_ _07045_ net563 vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__o211a_1
XANTENNA__12224__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17140_ clknet_leaf_81_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[5\]
+ _01369_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ net1258 vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__inv_2
XANTENNA__12775__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11564_ _07052_ _07051_ _07050_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__and3b_1
XFILLER_0_107_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11983__B1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09640__A2 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ net1082 team_04_WB.MEM_SIZE_REG_REG\[26\] team_04_WB.MEM_SIZE_REG_REG\[27\]
+ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__or3b_1
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17071_ clknet_leaf_48_wb_clk_i _00019_ _01300_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] net1095 net1053 vssd1 vssd1 vccd1
+ vccd1 _06082_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14283_ net1961 _03453_ _03455_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__a21oi_1
X_11495_ _05473_ _06980_ _06981_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or4b_1
XFILLER_0_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13724__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16022_ clknet_leaf_77_wb_clk_i _00005_ _00251_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09585__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10446_ _06023_ _06024_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__and2_1
X_13234_ net98 team_04_WB.MEM_SIZE_REG_REG\[7\] net984 vssd1 vssd1 vccd1 vccd1 _01669_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13724__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08826__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10377_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__inv_2
X_13165_ _07601_ net371 net290 net1767 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__a22o_1
XANTENNA__12305__A _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ net229 net678 vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__and2_1
X_13096_ _07528_ net367 net298 net1865 vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09156__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12047_ net232 net682 vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__and2_1
X_16924_ clknet_leaf_126_wb_clk_i _02593_ _01153_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15616__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14520__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08929__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09251__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08903__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16855_ clknet_leaf_174_wb_clk_i _02524_ _01084_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16786_ clknet_leaf_6_wb_clk_i _02455_ _01015_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13998_ _04972_ _03326_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15737_ net1296 vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__inv_2
X_12949_ net233 net2473 net320 vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XANTENNA__12463__A1 _06197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15668_ net1282 vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13007__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14619_ net1124 vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15599_ net1195 vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08140_ _03745_ _03750_ net730 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__mux2_1
XANTENNA__08514__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17338_ net1394 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__12766__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13963__A1 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__B1 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08071_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__mux2_1
Xclkload100 clknet_leaf_154_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload100/X sky130_fd_sc_hd__clkbuf_4
X_17269_ net1329 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
Xclkload111 clknet_leaf_160_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload111/X sky130_fd_sc_hd__clkbuf_4
Xclkload122 clknet_leaf_140_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload122/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_116_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12518__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload133 clknet_leaf_128_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__inv_6
Xclkload144 clknet_leaf_69_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload144/Y sky130_fd_sc_hd__inv_8
Xclkload155 clknet_leaf_97_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload155/X sky130_fd_sc_hd__clkbuf_8
Xclkload166 clknet_leaf_78_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload166/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_168_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload177 clknet_leaf_90_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload177/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12215__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _04558_ _04583_ net666 vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__mux2_2
XANTENNA__13745__S net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold17 net167 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ net1101 net1077 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__a21oi_1
Xhold28 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[20\]
+ vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\] vssd1 vssd1 vccd1
+ vccd1 net1476 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1009_A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09698__A2 _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11492__C _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _05130_ _05135_ net725 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1280_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout636_A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09456_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__mux2_1
XANTENNA__15969__Q team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08407_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09387_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1166_X net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08338_ net662 net660 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__X _07273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__mux2_1
XANTENNA__08830__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ _05895_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__inv_2
XANTENNA__12509__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ net576 _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08808__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _05561_ _05562_ _05646_ net621 _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__o311a_1
XFILLER_0_104_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13182__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__A0 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _05668_ _05772_ _05667_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_7_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__clkbuf_4
Xfanout1015 _06178_ vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08041__C net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 _03545_ vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10093_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] _04728_ vssd1
+ vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__or2_1
Xfanout1037 _03353_ vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__buf_2
X_14970_ net1151 vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1048 net1050 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12142__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\] vssd1 vssd1
+ vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_2
XANTENNA__13485__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ _03121_ _03144_ _03287_ _03243_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11496__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ clknet_leaf_137_wb_clk_i _02309_ _00869_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08992__S0 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13852_ _03516_ _07701_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__nand2_4
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _07327_ net2306 net323 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux2_1
X_16571_ clknet_leaf_97_wb_clk_i _02240_ _00800_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[544\]
+ sky130_fd_sc_hd__dfrtp_1
X_13783_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] net1044 _03173_
+ net1092 vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12445__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10995_ _06334_ _06336_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__a21bo_1
X_15522_ net1219 vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12734_ _07459_ net329 net400 net1771 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ net1155 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__inv_2
X_12665_ net246 net2530 net475 vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14404_ net1294 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__inv_2
XANTENNA__12748__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11616_ _05436_ _06248_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ net1205 vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12596_ _07565_ net480 net412 net2087 vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17123_ clknet_leaf_67_wb_clk_i _02758_ _01352_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14335_ net1190 vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
X_11547_ _06677_ _06886_ _07030_ _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__a22o_1
XANTENNA__09168__X _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17054_ clknet_leaf_50_wb_clk_i _00032_ _01283_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09609__A team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold509 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\] vssd1 vssd1
+ vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\] _03443_
+ net820 vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11858__B net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11478_ net571 _06807_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16005_ clknet_leaf_50_wb_clk_i _01681_ _00234_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_13217_ net85 team_04_WB.MEM_SIZE_REG_REG\[24\] net982 vssd1 vssd1 vccd1 vccd1 _01686_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13173__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] _06002_
+ _06003_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__o22ai_2
X_14197_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] _03404_
+ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[0\]
+ sky130_fd_sc_hd__and2b_1
XANTENNA__12035__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__C net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__A0 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12920__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ _07582_ net378 net296 net1965 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__a22o_1
XANTENNA__08800__X _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09129__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08659__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12133__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ net251 net2471 net302 vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__mux2_1
Xhold1209 team_04_WB.ADDR_START_VAL_REG\[0\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08337__C1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16907_ clknet_leaf_16_wb_clk_i _02576_ _01136_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\]
+ sky130_fd_sc_hd__dfrtp_1
X_16838_ clknet_leaf_20_wb_clk_i _02507_ _01067_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769_ clknet_leaf_135_wb_clk_i _02438_ _00998_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\]
+ sky130_fd_sc_hd__dfrtp_1
X_09310_ net628 _04919_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__or2_1
XANTENNA__12987__A2 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_752 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09241_ net727 _04851_ net712 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17259__1319 vssd1 vssd1 vccd1 vccd1 _17259__1319/HI net1319 sky130_fd_sc_hd__conb_1
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_90_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_118_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11114__A _06227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] net974 _04781_ vssd1 vssd1 vccd1
+ vccd1 _04783_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12739__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08123_ net721 _03733_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__nor2_1
XFILLER_0_160_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10953__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout217_A _07277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__mux2_1
XANTENNA__10982__A1_N _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap740 _03649_ vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
XANTENNA__13164__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12372__A0 _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12911__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07981__B team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08956_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__mux2_1
X_07907_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03522_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout753_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08887_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11883__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12427__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12819__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout639_X net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09508_ net725 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09701__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ net570 net555 net552 net533 vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__or4_4
XFILLER_0_149_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09439_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10566__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ net522 net603 _07455_ net429 net2311 vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_43_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11401_ _04724_ _04753_ net358 _06889_ net462 vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__o311a_1
XANTENNA__11959__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _07385_ net2509 net495 vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14335__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ team_04_WB.MEM_SIZE_REG_REG\[19\] net988 net981 team_04_WB.ADDR_START_VAL_REG\[19\]
+ net1005 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__o221a_1
XFILLER_0_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11332_ _06338_ _06482_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08333__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14051_ net5 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1
+ vccd1 vccd1 _01535_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_91_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11263_ net591 _04412_ net360 vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_162_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11166__A1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13002_ net603 _07462_ net471 net311 net1821 vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a32o_1
X_10214_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__and2b_1
XANTENNA__12902__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11194_ _06513_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__nand2_1
XANTENNA__11694__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _05698_ _05755_ _05699_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10076_ _04219_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] vssd1
+ vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__and2b_1
X_14953_ net1133 vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__inv_2
X_13904_ _02991_ _03278_ _02990_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08965__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14884_ net1189 vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__inv_2
X_16623_ clknet_leaf_187_wb_clk_i _02292_ _00852_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\]
+ sky130_fd_sc_hd__dfrtp_1
X_13835_ _02875_ _03225_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12418__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08098__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16554_ clknet_leaf_160_wb_clk_i _02223_ _00783_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\]
+ sky130_fd_sc_hd__dfrtp_1
X_13766_ team_04_WB.ADDR_START_VAL_REG\[19\] _03156_ vssd1 vssd1 vccd1 vccd1 _03157_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_139_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09295__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10978_ _04440_ _06465_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10757__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09103__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ net1272 vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__inv_2
XANTENNA__09390__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ net2145 net406 net343 _07409_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16485_ clknet_leaf_5_wb_clk_i _02154_ _00714_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\]
+ sky130_fd_sc_hd__dfrtp_1
X_13697_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15436_ net1122 vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__inv_2
X_12648_ _07619_ net488 net410 net1861 vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_84_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_154_Left_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ net1142 vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12579_ _07546_ net488 net418 net1660 vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17106_ clknet_leaf_63_wb_clk_i _02741_ _01335_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14318_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_113_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold306 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\] vssd1 vssd1
+ vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
X_15298_ net1218 vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__inv_2
Xhold317 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\] vssd1 vssd1
+ vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\] vssd1 vssd1
+ vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ clknet_leaf_41_wb_clk_i _02706_ _01266_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold339 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\] vssd1 vssd1
+ vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13146__A2 net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14249_ _03433_ _03434_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11157__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout808 _03550_ vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__clkbuf_4
Xfanout819 net821 vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10904__A1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08810_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__mux2_1
XANTENNA__08389__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09790_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__mux2_1
Xhold1006 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\] vssd1 vssd1
+ vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_163_Left_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1017 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\] vssd1 vssd1
+ vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\]
+ net870 vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
Xhold1028 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[2\] vssd1
+ vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13854__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\] vssd1 vssd1
+ vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10668__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09361__X _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12409__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09013__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout334_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13909__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_172_Left_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__mux2_1
XANTENNA__13978__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09155_ _04762_ _04763_ _04764_ _04765_ net788 net809 vssd1 vssd1 vccd1 vccd1 _04766_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12374__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout501_A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12227__X _07556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1243_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12593__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09086_ _03634_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13137__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13994__A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08037_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net974 _03647_ vssd1 vssd1 vccd1
+ vccd1 _03648_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold840 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\] vssd1 vssd1
+ vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\] vssd1 vssd1
+ vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\] vssd1 vssd1
+ vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold873 _02721_ vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\] vssd1 vssd1
+ vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15982__Q team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold895 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\] vssd1 vssd1
+ vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout968_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14098__B1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ net626 _05058_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nand2_1
XANTENNA__08299__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_157_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08939_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__mux2_1
XANTENNA__13845__B1 _03235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Right_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__A team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15714__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11950_ net691 _07410_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10901_ _05056_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__nor2_1
XANTENNA__09712__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07354_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_28_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12549__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13620_ _07039_ net271 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__nand2_1
X_10832_ net644 _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11084__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13551_ _02934_ _02940_ team_04_WB.ADDR_START_VAL_REG\[20\] vssd1 vssd1 vccd1 vccd1
+ _02942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10763_ net466 _06250_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ _07499_ net493 net427 net2039 vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a22o_1
X_16270_ clknet_leaf_32_wb_clk_i _01939_ _00499_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[243\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14022__B1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ team_04_WB.ADDR_START_VAL_REG\[28\] _02865_ _02869_ _02872_ vssd1 vssd1 vccd1
+ vccd1 _02873_ sky130_fd_sc_hd__and4_1
XANTENNA_input97_A wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _05280_ _06181_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ net1208 vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12433_ net2103 net434 _07637_ net524 vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XANTENNA__10593__A team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11387__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ net1160 vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12364_ net217 net2457 net496 vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17149__Q team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14103_ team_04_WB.MEM_SIZE_REG_REG\[2\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[2\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_168_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11315_ net572 _06803_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nand2_1
XANTENNA__13128__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15083_ net1160 vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12295_ net211 net669 vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__and2_1
XANTENNA__09593__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14034_ net23 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1
+ vccd1 vccd1 _01552_ sky130_fd_sc_hd__o22a_1
XANTENNA__09201__B1 _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246_ net559 _06664_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__or2_1
XANTENNA__10532__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ net553 _06663_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17258__1318 vssd1 vssd1 vccd1 vccd1 _17258__1318/HI net1318 sky130_fd_sc_hd__conb_1
X_10128_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _05342_ _05737_
+ _05735_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__a31o_1
XANTENNA__12639__A1 _07610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15985_ clknet_leaf_52_wb_clk_i _01661_ _00214_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08938__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _03894_ vssd1
+ vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__and2_1
X_14936_ net1222 vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_106_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14867_ net1237 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ team_04_WB.ADDR_START_VAL_REG\[25\] _03201_ _03205_ _03208_ vssd1 vssd1 vccd1
+ vccd1 _03209_ sky130_fd_sc_hd__and4_1
X_16606_ clknet_leaf_129_wb_clk_i _02275_ _00835_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\]
+ sky130_fd_sc_hd__dfrtp_1
X_14798_ net1200 vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16537_ clknet_leaf_178_wb_clk_i _02206_ _00766_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13749_ team_04_WB.ADDR_START_VAL_REG\[8\] _03139_ vssd1 vssd1 vccd1 vccd1 _03140_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_35_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10822__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16468_ clknet_leaf_8_wb_clk_i _02137_ _00697_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15419_ net1136 vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16399_ clknet_leaf_184_wb_clk_i _02068_ _00628_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_171_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12575__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[8\] vssd1 vssd1
+ vccd1 vccd1 net1540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12207__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold114 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[2\]
+ vssd1 vssd1 vccd1 vccd1 net1551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13119__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[26\]
+ vssd1 vssd1 vccd1 vccd1 net1562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[28\] vssd1
+ vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14703__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold147 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\] vssd1 vssd1
+ vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\] vssd1 vssd1
+ vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _03612_ _03637_ _05443_ _05521_ net759 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__a41o_1
Xhold169 _02720_ vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout605 net606 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__buf_2
Xfanout616 _06192_ vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09445__A1_N net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09743__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _03893_ _03947_ _04002_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nor4_1
Xfanout627 _04947_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
Xfanout638 _04273_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_2
Xfanout649 _07520_ vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__buf_4
XANTENNA__10353__A2 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09773_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08724_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\]
+ net904 vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__mux2_1
XANTENNA__13968__A_N _04192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ _04262_ _04263_ _04264_ _04265_ net783 net805 vssd1 vssd1 vccd1 vccd1 _04266_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12369__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08586_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09354__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08582__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12566__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09138_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12030__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11796__X _07280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11021__B team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09069_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__mux2_1
X_11100_ _06588_ _06247_ _06240_ _06578_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ net237 net676 vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__and2_2
XANTENNA__08170__X _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\] vssd1 vssd1
+ vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold681 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\] vssd1 vssd1
+ vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold692 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\] vssd1 vssd1
+ vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ _06499_ _06519_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15444__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ net1289 vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_86_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08757__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ _07634_ net472 net316 net2080 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XANTENNA__12097__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input12_A DAT_I[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ net1148 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__inv_2
X_11933_ net688 _06200_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__and2_2
XANTENNA__11844__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14652_ net1126 vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__inv_2
X_11864_ net694 _06781_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13603_ _02981_ _02990_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__nand2_1
X_10815_ _06282_ _06300_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__nand3_2
X_14583_ net1179 vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11795_ net757 _05815_ _06185_ net660 net689 vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_60_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ clknet_leaf_145_wb_clk_i _01991_ _00551_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09588__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _07843_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07897__A team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08607__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10746_ net639 net549 _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08473__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_147_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_147_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16253_ clknet_leaf_131_wb_clk_i _01922_ _00482_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\]
+ sky130_fd_sc_hd__dfrtp_1
X_13465_ _06625_ net272 net709 vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10677_ net2667 net1017 net1013 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1
+ vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
XANTENNA__08064__Y _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15204_ net1189 vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__inv_2
XANTENNA__12557__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08225__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ net521 net605 _07350_ net433 net1624 vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a32o_1
X_16184_ clknet_leaf_153_wb_clk_i _01853_ _00413_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\]
+ sky130_fd_sc_hd__dfrtp_1
X_13396_ _07758_ _07821_ _07757_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12027__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10032__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput208 net208 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
X_15135_ net1250 vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__inv_2
XANTENNA__08320__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ net223 net670 vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__and2_1
XANTENNA__14523__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ net1151 vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__inv_2
XANTENNA__11866__B net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ net233 net674 vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__and2_1
X_14017_ net1537 net1073 _03344_ net265 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a22o_1
X_11229_ net575 _06642_ _06717_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12043__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10335__A2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__C1 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ clknet_leaf_51_wb_clk_i _01644_ _00197_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_125_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14919_ net1134 vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__inv_2
X_15899_ clknet_leaf_35_wb_clk_i _01576_ _00126_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08440_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[760\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08139__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08371_ _03978_ _03979_ _03980_ _03981_ net784 net808 vssd1 vssd1 vccd1 vccd1 _03982_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12796__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09498__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13321__B team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12012__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_X clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1039_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09527__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout402 _07669_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_6
XANTENNA_fanout499_A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 net415 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
XANTENNA__08075__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout424 _07656_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1206_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout435 _07625_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12720__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 net449 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input4_A DAT_I[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net461 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_4
X_09825_ _05404_ net541 vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__xnor2_1
Xfanout468 net469 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout666_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 net480 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout287_X net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ net726 _05366_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or2_1
XANTENNA__12079__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\]
+ net937 vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11826__A2 _07305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout833_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12400__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08638_ _04218_ _04245_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ net728 _04179_ net712 vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10600_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[0\]
+ _06138_ net1049 vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__mux2_1
XANTENNA__12787__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11580_ _06268_ _06615_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12251__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[23\]
+ _06092_ net1047 vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257__1317 vssd1 vssd1 vccd1 vccd1 _17257__1317/HI net1317 sky130_fd_sc_hd__conb_1
XFILLER_0_162_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ net87 team_04_WB.ADDR_START_VAL_REG\[26\] net975 vssd1 vssd1 vccd1 vccd1
+ _01656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _06030_
+ _06035_ _06040_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a311o_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12201_ net254 net647 vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _07617_ net378 net292 net1672 vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a22o_1
X_10393_ net279 _05976_ _05977_ _05973_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07966__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ net227 net2534 net512 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10590__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ net1904 net354 _07486_ net450 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a22o_1
X_16940_ clknet_leaf_112_wb_clk_i _02609_ _01169_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09802__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ team_04_WB.MEM_SIZE_REG_REG\[8\] _06502_ vssd1 vssd1 vccd1 vccd1 _06503_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16871_ clknet_leaf_165_wb_clk_i _02540_ _01100_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout980 net981 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__buf_4
Xfanout991 _07692_ vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_4
X_15822_ clknet_leaf_93_wb_clk_i _01499_ _00049_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11278__A0 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15753_ net1267 vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__inv_2
XANTENNA__09566__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13406__B team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _07631_ net469 net314 net1716 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ net688 _07382_ _07383_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__a21bo_1
X_14704_ net1165 vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15684_ net1268 vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ _07598_ net327 net384 net2054 vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__a22o_1
X_14635_ net1161 vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11847_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net269 vssd1 vssd1 vccd1 vccd1
+ _07324_ sky130_fd_sc_hd__and2_1
XANTENNA__14518__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12778__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14566_ net1185 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11778_ net653 net214 vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09111__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A0 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ team_04_WB.ADDR_START_VAL_REG\[23\] _02901_ _02907_ vssd1 vssd1 vccd1 vccd1
+ _02908_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16305_ clknet_leaf_180_wb_clk_i _01974_ _00534_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\]
+ sky130_fd_sc_hd__dfrtp_1
X_17285_ net1341 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10729_ net628 net627 net552 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__mux2_1
X_14497_ net1164 vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16236_ clknet_4_12__leaf_wb_clk_i _01905_ _00465_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\]
+ sky130_fd_sc_hd__dfrtp_1
X_13448_ _07727_ _07873_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__nand2_1
Xclkload12 clknet_leaf_186_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_6
Xclkload23 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__08950__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload34 clknet_leaf_179_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload34/X sky130_fd_sc_hd__clkbuf_8
Xclkload45 clknet_leaf_166_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload45/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__13742__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16167_ clknet_leaf_24_wb_clk_i _01836_ _00396_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload56 clknet_leaf_33_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_2
X_13379_ _07770_ _07771_ _07772_ _07804_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__o22a_1
Xclkload67 clknet_leaf_48_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload67/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10781__A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload78 clknet_leaf_40_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload78/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11753__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12950__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_149_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15118_ net1197 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__inv_2
Xclkload89 clknet_leaf_143_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_149_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16098_ clknet_leaf_145_wb_clk_i _01767_ _00327_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07940_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net973 _03549_ vssd1 vssd1 vccd1
+ vccd1 _03551_ sky130_fd_sc_hd__o21ai_2
X_15049_ net1132 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_44_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12702__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09610_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\] net1010
+ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13258__A1 team_04_WB.ADDR_START_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__X _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08397__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ _05148_ _05149_ _05150_ _05151_ net793 net802 vssd1 vssd1 vccd1 vccd1 _05152_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11808__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09472_ _05065_ _05071_ _05082_ net718 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a22o_4
XFILLER_0_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12481__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12769__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_A _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13332__A team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08354_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\]
+ net862 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12233__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08426__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09021__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10244__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_8
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08285_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__mux2_1
XANTENNA__13981__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout414_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09528__Y _05139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12941__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout783_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1209 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
Xfanout221 net222 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout1219 net1220 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09691__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout232 _07420_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_2
Xfanout243 _07374_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
XANTENNA_fanout950_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 _07380_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _05415_ _05416_ _05417_ _05418_ net834 net738 vssd1 vssd1 vccd1 vccd1 _05419_
+ sky130_fd_sc_hd__mux4_1
Xfanout287 _06205_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__buf_4
XANTENNA__13249__A1 team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _07682_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13523__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09548__S0 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08100__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10569__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12750_ _07475_ net342 net402 net2011 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08676__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12472__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11701_ net572 _07189_ _07188_ net582 vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__a211o_1
XFILLER_0_167_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08771__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ net231 net2506 net477 vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__mux2_1
XANTENNA__14338__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14420_ net1267 vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11632_ net466 _06808_ _06809_ _06884_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o211a_1
XANTENNA__12224__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09625__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11432__A0 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14351_ net1191 vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ net565 _05475_ _06273_ _06248_ _05380_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13302_ net1082 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 _07728_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11983__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17070_ clknet_leaf_48_wb_clk_i _00017_ _01299_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10514_ _06081_ net1582 net1022 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
Xwire644 _03780_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14282_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[22\] _03453_
+ net821 vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_98_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08770__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ _04923_ net365 net358 _04921_ _06982_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__o221a_1
X_16021_ clknet_leaf_78_wb_clk_i _00004_ _00250_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13185__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ net99 team_04_WB.MEM_SIZE_REG_REG\[8\] net984 vssd1 vssd1 vccd1 vccd1 _01670_
+ sky130_fd_sc_hd__mux2_1
X_10445_ _06016_ _06021_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12932__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _07600_ net369 net290 net1848 vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10376_ _05962_ _05959_ net282 vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12305__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ net2542 net354 _07512_ net451 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13095_ _07527_ net374 net299 net1847 vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12046_ net2357 net517 _07476_ net454 vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a22o_1
XANTENNA__11499__B1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16923_ clknet_leaf_97_wb_clk_i _02592_ _01152_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10540__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12321__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16854_ clknet_leaf_12_wb_clk_i _02523_ _01083_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09106__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16785_ clknet_leaf_172_wb_clk_i _02454_ _01014_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\]
+ sky130_fd_sc_hd__dfrtp_1
X_13997_ net1454 net1065 _03333_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12999__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15736_ net1295 vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__inv_2
X_12948_ net261 net2439 net320 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12463__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_162_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_162_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15667_ net1284 vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__inv_2
X_12879_ _07579_ net330 net388 net2079 vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14618_ net1146 vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15598_ net1197 vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17337_ net1393 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
X_14549_ net1178 vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__inv_2
XANTENNA__09711__S0 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08514__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13963__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11423__B1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09776__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ net728 _03680_ net713 vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__o21a_1
XANTENNA__08680__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17268_ net1328 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xclkload101 clknet_leaf_155_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload101/X sky130_fd_sc_hd__clkbuf_8
Xclkload112 clknet_leaf_162_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_116_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload123 clknet_leaf_141_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__bufinv_16
Xclkload134 clknet_leaf_63_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload134/Y sky130_fd_sc_hd__inv_6
XANTENNA__13176__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload145 clknet_leaf_70_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload145/Y sky130_fd_sc_hd__inv_6
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16219_ clknet_leaf_101_wb_clk_i _01888_ _00448_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\]
+ sky130_fd_sc_hd__dfrtp_1
X_17199_ clknet_leaf_59_wb_clk_i _02811_ _01428_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload156 clknet_leaf_98_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload156/Y sky130_fd_sc_hd__bufinv_16
Xclkload167 clknet_leaf_80_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload167/Y sky130_fd_sc_hd__inv_8
XANTENNA__12923__A0 _07246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_168_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload178 clknet_leaf_94_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload178/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_12_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12215__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12930__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ net718 _04582_ _04571_ _04570_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__13479__A1 _05800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ _03535_ _03536_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__and2_1
XANTENNA_wire637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\] vssd1 vssd1
+ vccd1 vccd1 net1455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\] vssd1 vssd1 vccd1
+ vccd1 net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17256__1316 vssd1 vssd1 vccd1 vccd1 _17256__1316/HI net1316 sky130_fd_sc_hd__conb_1
XFILLER_0_78_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17238__1404 vssd1 vssd1 vccd1 vccd1 net1404 _17238__1404/LO sky130_fd_sc_hd__conb_1
XANTENNA__09016__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout364_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _05131_ _05132_ _05133_ _05134_ net832 net747 vssd1 vssd1 vccd1 vccd1 _05135_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08855__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08753__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout531_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_A _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1273_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08406_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__mux2_1
X_09386_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__mux2_1
XANTENNA__12206__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08337_ _03639_ _03641_ _03947_ net752 _03725_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a221oi_2
XANTENNA__14308__D net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11965__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07995__A team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08830__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08268_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux2_1
XANTENNA__08830__B2 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout998_A _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ net644 _03808_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12406__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12914__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ _05561_ _05562_ _05646_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14116__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _05670_ _05672_ _05770_ _05671_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_7_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 _06154_ vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__clkbuf_4
Xfanout1016 net1018 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_58_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08041__D net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14131__A2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1027 _03545_ vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10092_ _05700_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor2_1
Xfanout1038 _03352_ vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_2
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1049 net1050 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__buf_4
XANTENNA__09543__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ net1040 _03289_ _03290_ net1071 net1495 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a32o_1
XANTENNA__12693__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__A3 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13851_ _02853_ _03231_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08992__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _07320_ net2497 net322 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__mux2_1
XANTENNA__11980__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13782_ _07825_ _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
X_16570_ clknet_leaf_36_wb_clk_i _02239_ _00799_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ net641 _06333_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_48_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _07458_ net327 net400 net2157 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15521_ net1129 vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__inv_2
XANTENNA__12996__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__A team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15452_ net1145 vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_67_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12664_ net236 net2511 net475 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14403_ net1289 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11405__A0 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11979__X _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11615_ _05379_ _06412_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__xnor2_1
X_15383_ net1233 vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12595_ _07564_ net481 net412 net2015 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11956__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334_ net1191 vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__inv_2
X_17122_ clknet_leaf_63_wb_clk_i _02757_ _01351_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11546_ net576 _07031_ _06278_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13158__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17053_ clknet_leaf_47_wb_clk_i _00029_ _01282_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14265_ _03443_ _03444_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10535__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _06959_ _06965_ net585 vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16004_ clknet_leaf_50_wb_clk_i _01680_ _00233_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11220__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13216_ net86 team_04_WB.MEM_SIZE_REG_REG\[25\] net983 vssd1 vssd1 vccd1 vccd1 _01687_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12905__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] _06006_
+ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_164_Right_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14196_ _03403_ _03366_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12035__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14107__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13846__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _07581_ net379 net296 net1871 vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a22o_1
X_10359_ _05944_ _05947_ net618 vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10392__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14122__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13078_ net253 net2330 net302 vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__mux2_1
X_16906_ clknet_leaf_162_wb_clk_i _02575_ _01135_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\]
+ sky130_fd_sc_hd__dfrtp_1
X_12029_ _07368_ net684 vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__and2_1
XANTENNA__09168__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16837_ clknet_leaf_185_wb_clk_i _02506_ _01066_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11892__B1 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16768_ clknet_leaf_140_wb_clk_i _02437_ _00997_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13633__B2 net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15719_ net1294 vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16699_ clknet_leaf_100_wb_clk_i _02368_ _00928_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\]
+ sky130_fd_sc_hd__dfrtp_1
X_09240_ _04847_ _04848_ _04849_ _04850_ net824 net733 vssd1 vssd1 vccd1 vccd1 _04851_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13936__A2 net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] net974 _04781_ vssd1 vssd1 vccd1
+ vccd1 _04782_ sky130_fd_sc_hd__o21a_2
XFILLER_0_111_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12925__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14706__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11947__A1 net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11947__B2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ _03729_ _03730_ _03731_ _03732_ net825 net750 vssd1 vssd1 vccd1 vccd1 _03733_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13149__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08053_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12226__A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11175__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10383__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A _06073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14113__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__B _07165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout481_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__inv_2
X_08886_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12427__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09507_ _05114_ _05115_ _05116_ _05117_ net832 net737 vssd1 vssd1 vccd1 vccd1 _05118_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12978__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _05045_ _05046_ _05047_ _05048_ net793 net813 vssd1 vssd1 vccd1 vccd1 _05049_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13520__A _06681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_391 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11400_ _04724_ _04753_ net361 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11959__B net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _07380_ net2450 net495 vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08614__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11331_ _06514_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_158_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ net6 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1
+ vccd1 vccd1 _01536_ sky130_fd_sc_hd__o22a_1
XFILLER_0_162_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11262_ net566 _06741_ _06739_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_91_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11166__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ net600 _07461_ net468 net310 net1885 vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a32o_1
XFILLER_0_162_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13560__B1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _05768_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__xor2_1
X_11193_ team_04_WB.MEM_SIZE_REG_REG\[22\] _06512_ vssd1 vssd1 vccd1 vccd1 _06682_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__14351__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10913__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14104__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__B _07182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _05702_ _05754_ _05701_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12115__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _04274_ vssd1
+ vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__and2_1
X_14952_ net1117 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__inv_2
X_13903_ _03098_ _03143_ _03145_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__o21a_1
XANTENNA__10677__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11874__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08965__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14883_ net1175 vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__inv_2
X_16622_ clknet_leaf_26_wb_clk_i _02291_ _00851_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\]
+ sky130_fd_sc_hd__dfrtp_1
X_13834_ _03222_ _03224_ _02900_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__o21a_1
XFILLER_0_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12418__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ net997 _03152_ _03155_ _03149_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__o211a_1
X_16553_ clknet_leaf_123_wb_clk_i _02222_ _00782_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__B1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12969__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ _04440_ _06465_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__or2_1
XANTENNA__09295__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13091__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15504_ net1166 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12716_ net2115 net406 net343 _07403_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a22o_1
X_13696_ _03045_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09390__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16484_ clknet_leaf_168_wb_clk_i _02153_ _00713_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[457\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12647_ _07618_ net490 net410 net1632 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
X_15435_ net1122 vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14526__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14040__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11929__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15366_ net1110 vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__inv_2
X_12578_ _07545_ net492 net419 net1987 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a22o_1
X_17255__1315 vssd1 vssd1 vccd1 vccd1 _17255__1315/HI net1315 sky130_fd_sc_hd__conb_1
X_17105_ clknet_leaf_63_wb_clk_i _02740_ _01334_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14317_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[23\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[22\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[19\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[18\] net1091
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\] vssd1 vssd1
+ vccd1 vccd1 _03477_ sky130_fd_sc_hd__mux4_1
X_17237__1403 vssd1 vssd1 vccd1 vccd1 net1403 _17237__1403/LO sky130_fd_sc_hd__conb_1
X_11529_ _05003_ _05030_ net361 vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_152_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15297_ net1167 vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__inv_2
Xhold307 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\] vssd1 vssd1
+ vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 net127 vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] _03432_ net820
+ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o21ai_1
Xhold329 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\] vssd1 vssd1
+ vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ clknet_leaf_112_wb_clk_i _02705_ _01265_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12354__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ _03514_ _03392_ _03378_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12333__X _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net811 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10904__A2 _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08740_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\]
+ net870 vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
Xhold1007 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\] vssd1 vssd1
+ vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\] vssd1 vssd1
+ vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\] vssd1 vssd1
+ vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10668__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08671_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12409__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12655__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1069_A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09154_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08105_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09085_ net703 _04669_ _04386_ net666 vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1236_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08036_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[22\] net1009
+ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput90 wbs_dat_i[29] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_1
XANTENNA__13994__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold830 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\] vssd1 vssd1
+ vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold841 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\] vssd1 vssd1
+ vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout696_A _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold852 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\] vssd1 vssd1
+ vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold863 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1011\] vssd1 vssd1
+ vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12390__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\] vssd1 vssd1
+ vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\] vssd1 vssd1
+ vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\] vssd1 vssd1
+ vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_09987_ _05056_ _05058_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout863_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ _04545_ _04546_ _04547_ _04548_ net792 net812 vssd1 vssd1 vccd1 vccd1 _04549_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12648__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13845__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12122__C net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__B team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_X net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10900_ _05084_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__xnor2_1
X_11880_ _05468_ _06200_ _07216_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__and3_2
XFILLER_0_93_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09204__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10831_ _03808_ _06309_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ team_04_WB.ADDR_START_VAL_REG\[20\] _02934_ _02940_ vssd1 vssd1 vccd1 vccd1
+ _02941_ sky130_fd_sc_hd__and3_1
XANTENNA__11084__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10762_ _05447_ _05470_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11623__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12501_ _07498_ net483 net425 net1724 vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a22o_1
XANTENNA__08047__C net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13783__A2_N net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ net997 _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10693_ _05280_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14346__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15220_ net1227 vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12432_ net653 net608 net229 vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10593__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15151_ net1196 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12363_ net219 net2405 net495 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14102_ team_04_WB.MEM_SIZE_REG_REG\[1\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[1\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__o221a_2
XANTENNA__11792__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11314_ _06801_ _06802_ net559 vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15082_ net1105 vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__inv_2
X_12294_ _05221_ _06194_ _07590_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__or3_4
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ net25 net1062 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1
+ vccd1 vccd1 _01553_ sky130_fd_sc_hd__a22o_1
XANTENNA__12336__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ _06711_ _06733_ net463 vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09201__B2 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12887__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11176_ net553 _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nor2_1
XANTENNA__12313__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08960__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__X _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _05735_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__and2b_1
X_15984_ clknet_leaf_52_wb_clk_i _01660_ _00213_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12639__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10058_ _05667_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__and2b_1
X_14935_ net1231 vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__inv_2
XANTENNA__08938__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14866_ net1238 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09114__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16605_ clknet_leaf_132_wb_clk_i _02274_ _00834_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\]
+ sky130_fd_sc_hd__dfrtp_1
X_13817_ net1002 _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_158_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14797_ net1210 vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_69_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11075__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16536_ clknet_leaf_151_wb_clk_i _02205_ _00765_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\]
+ sky130_fd_sc_hd__dfrtp_1
X_13748_ net999 _03135_ _03138_ _03133_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16467_ clknet_leaf_182_wb_clk_i _02136_ _00696_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ team_04_WB.MEM_SIZE_REG_REG\[1\] net993 net991 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ net1000 vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_14_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15418_ net1142 vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__inv_2
X_16398_ clknet_leaf_26_wb_clk_i _02067_ _00627_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08254__A _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15349_ net1207 vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__inv_2
Xhold104 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[7\] vssd1
+ vssd1 vccd1 vccd1 net1541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09784__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold115 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[17\] vssd1
+ vssd1 vccd1 vccd1 net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09637__X _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[15\]
+ vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold137 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[12\]
+ vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold148 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[15\] vssd1
+ vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09910_ _05464_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold159 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\] vssd1 vssd1
+ vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15087__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17019_ clknet_leaf_97_wb_clk_i _02688_ _01248_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12878__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net612 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__buf_2
X_09841_ _03644_ _03727_ _03782_ _03835_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or4_1
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__buf_2
Xfanout628 _04892_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12223__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout639 _04218_ vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09772_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__mux2_1
X_08723_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\]
+ net870 vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_13_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout277_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08654_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09024__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08585_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout444_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09354__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12385__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09206_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09137_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09068_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\]
+ net873 vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout980_A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08019_ _03598_ _03617_ _03620_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__or3_4
XANTENNA__12318__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold660 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\] vssd1 vssd1
+ vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12869__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold671 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\] vssd1 vssd1
+ vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11030_ team_04_WB.MEM_SIZE_REG_REG\[31\] _06518_ vssd1 vssd1 vccd1 vccd1 _06519_
+ sky130_fd_sc_hd__xor2_1
Xhold682 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\] vssd1 vssd1
+ vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\] vssd1 vssd1
+ vccd1 vccd1 net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ net608 _07403_ net472 net316 net1545 vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a32o_1
XANTENNA__11829__B1 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17254__1314 vssd1 vssd1 vccd1 vccd1 _17254__1314/HI net1314 sky130_fd_sc_hd__conb_1
X_14720_ net1213 vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__inv_2
X_11932_ net1968 net529 net458 _07397_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a22o_1
X_17236__1402 vssd1 vssd1 vccd1 vccd1 net1402 _17236__1402/LO sky130_fd_sc_hd__conb_1
XANTENNA__08170__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11863_ net688 _07337_ _07336_ _07335_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__a211o_1
X_14651_ net1124 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13046__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ _02970_ _02992_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ _04140_ _04193_ _05463_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ net1185 vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__inv_2
X_11794_ net2167 net527 net445 _07278_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16321_ clknet_leaf_141_wb_clk_i _01990_ _00550_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13533_ _07837_ _07840_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ net638 net543 vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and2_1
XANTENNA__08473__A2 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13464_ _02853_ _02854_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__nand2_1
X_16252_ clknet_leaf_127_wb_clk_i _01921_ _00481_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ net1599 net1018 net1014 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1
+ vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15203_ net1170 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__inv_2
X_12415_ net525 net610 _07341_ net435 net1550 vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a32o_1
XANTENNA__11987__X _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _07763_ _07820_ _07762_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16183_ clknet_leaf_161_wb_clk_i _01852_ _00412_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12346_ net2500 net501 _07617_ net453 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
X_15134_ net1215 vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__inv_2
Xoutput209 net209 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_187_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_187_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__07984__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15065_ net1248 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__inv_2
XANTENNA__10543__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net2460 net505 _07581_ net453 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
XANTENNA__11517__C1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09109__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ _05374_ _03336_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__nor2_1
X_11228_ net571 _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__nand2_1
XANTENNA__12043__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11159_ _06227_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_108_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15967_ clknet_leaf_47_wb_clk_i _01643_ _00196_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_125_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14918_ net1105 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15898_ clknet_leaf_99_wb_clk_i _01575_ _00125_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14849_ net1130 vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__inv_2
XANTENNA__13037__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09779__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[441\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__mux2_1
XANTENNA__08683__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_173_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16519_ clknet_leaf_24_wb_clk_i _02188_ _00748_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13993__B1 _03331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12548__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11897__X _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12933__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09019__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout403 _07669_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_2
Xfanout414 net415 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08075__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout425 _07656_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__clkbuf_4
Xfanout436 net444 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_4
XANTENNA_fanout394_A _07672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
X_09824_ net661 _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout1101_A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__clkbuf_4
Xfanout469 _07668_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_14__f_wb_clk_i clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09755_ _05362_ _05363_ _05364_ _05365_ net837 net739 vssd1 vssd1 vccd1 vccd1 _05366_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout561_A _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\]
+ net937 vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
X_09686_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08637_ net639 _04245_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1091_X net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13028__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08568_ _04175_ _04176_ _04177_ _04178_ net825 net734 vssd1 vssd1 vccd1 vccd1 _04179_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10695__Y _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_30_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout614_X net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08499_ _04106_ _04107_ _04108_ _04109_ net784 net808 vssd1 vssd1 vccd1 vccd1 _04110_
+ sky130_fd_sc_hd__mux4_1
X_10530_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net1095 net1052 vssd1 vssd1 vccd1
+ vccd1 _06092_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12539__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _06036_
+ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14624__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ net2518 net508 _07541_ net449 vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a22o_1
XANTENNA__11600__X _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _07616_ net377 net292 net2058 vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10392_ _05619_ net624 _05971_ net283 vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07966__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ net217 net2447 net512 vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10590__C net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12062_ net213 net678 vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__and2_2
XFILLER_0_25_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold490 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\] vssd1 vssd1
+ vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ team_04_WB.MEM_SIZE_REG_REG\[7\] team_04_WB.MEM_SIZE_REG_REG\[6\] _06501_
+ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_53_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ clknet_leaf_20_wb_clk_i _02539_ _01099_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08768__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__clkbuf_2
Xfanout981 _07707_ vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__buf_4
X_15821_ clknet_leaf_84_wb_clk_i _01498_ _00048_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout992 _07690_ vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10599__A team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11278__A1 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15752_ net1269 vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__inv_2
XANTENNA__09566__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ _07630_ net468 net314 net1587 vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1190 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\] vssd1 vssd1
+ vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_103_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ net1140 vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__inv_2
X_11915_ _03632_ _05937_ _05941_ net756 net691 vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__o221a_1
X_15683_ net1268 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12895_ _07597_ net334 net385 net1788 vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__a22o_1
XANTENNA_output209_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09599__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ net1124 vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__inv_2
X_11846_ net704 _05867_ _07322_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12778__A1 _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_166_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14565_ net1184 vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__inv_2
XANTENNA__10538__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ _06186_ _06624_ _07263_ net615 vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__a211oi_2
XANTENNA__08446__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16304_ clknet_leaf_1_wb_clk_i _01973_ _00533_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\]
+ sky130_fd_sc_hd__dfrtp_1
X_13516_ _02904_ _02906_ net996 vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__mux2_1
XANTENNA__11450__A1 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ _06213_ _06216_ net563 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__mux2_1
X_17284_ net1340 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_83_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14496_ net1251 vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16235_ clknet_leaf_22_wb_clk_i _01904_ _00464_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\]
+ sky130_fd_sc_hd__dfrtp_1
X_13447_ _07871_ _07872_ _07726_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__o21bai_1
X_10659_ net1575 net1017 net1013 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1
+ vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload13 clknet_leaf_187_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__inv_6
Xclkload24 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_70_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload35 clknet_leaf_180_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload35/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_125_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload46 clknet_leaf_168_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__bufinv_16
X_13378_ _07776_ _07803_ _07775_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__o21ba_1
X_16166_ clknet_leaf_18_wb_clk_i _01835_ _00395_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload57 clknet_leaf_34_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__inv_8
XANTENNA__10781__B net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload68 clknet_leaf_49_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_6
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload79 clknet_leaf_41_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload79/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_77_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15117_ net1152 vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12329_ net256 net671 vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_149_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16097_ clknet_leaf_136_wb_clk_i _01766_ _00326_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15048_ net1118 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_166_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08678__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16999_ clknet_leaf_165_wb_clk_i _02668_ _01228_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09540_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\]
+ net951 vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__mux2_1
XANTENNA__12466__B1 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09471_ _05076_ _05081_ net724 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__mux2_1
XANTENNA__12928__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08422_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__mux2_1
XANTENNA__13613__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10956__B _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09302__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\]
+ net862 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08284_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload7 clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13981__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12663__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10972__A _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1051_A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A _07664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17253__1313 vssd1 vssd1 vccd1 vccd1 _17253__1313/HI net1313 sky130_fd_sc_hd__conb_1
XFILLER_0_30_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17235__1401 vssd1 vssd1 vccd1 vccd1 net1401 _17235__1401/LO sky130_fd_sc_hd__conb_1
XFILLER_0_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10401__C1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08070__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout211 _07246_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1209 net1254 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__buf_2
XANTENNA_fanout776_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 _07432_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 net235 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
Xfanout244 _07340_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_2
XFILLER_0_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout255 _07368_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 _07234_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__buf_4
XFILLER_0_5_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout277 net279 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
X_09807_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1\]
+ net890 vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__mux2_1
Xfanout288 _06526_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
X_07999_ team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] net1080 net1029 net1025 vssd1
+ vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__and4_1
Xfanout299 _07682_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout943_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Left_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09548__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ net748 _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__nor2_1
X_15804__23 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__inv_2
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] net974 _05278_ vssd1 vssd1 vccd1
+ vccd1 _05280_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11700_ _06553_ _06560_ net559 vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__mux2_1
X_12680_ net223 net2561 net477 vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09212__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13957__B1 _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ _06418_ _06420_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_64_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09625__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14350_ net1191 vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_145_Right_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11432__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ _05336_ net548 net358 vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13301_ team_04_WB.MEM_SIZE_REG_REG\[29\] _07726_ vssd1 vssd1 vccd1 vccd1 _07727_
+ sky130_fd_sc_hd__nand2_1
X_10513_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[29\]
+ _06080_ net1047 vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11983__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14281_ _03453_ _03454_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__nor2_1
XANTENNA__10882__A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11493_ _04922_ net362 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__nand2_1
XANTENNA__14354__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13232_ net100 team_04_WB.MEM_SIZE_REG_REG\[9\] net984 vssd1 vssd1 vccd1 vccd1 _01671_
+ sky130_fd_sc_hd__mux2_1
X_16020_ clknet_leaf_77_wb_clk_i _00003_ _00249_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_10444_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _06022_
+ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09448__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input72_A wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07939__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _07599_ net368 net290 net1986 vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10375_ _05621_ _05960_ _05961_ net624 vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ net231 net678 vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13094_ _07526_ net369 net299 net1770 vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16922_ clknet_leaf_38_wb_clk_i _02591_ _01151_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ net223 net683 vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12696__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16853_ clknet_leaf_12_wb_clk_i _02522_ _01082_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12321__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_161_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10122__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16784_ clknet_leaf_190_wb_clk_i _02453_ _01013_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08116__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13996_ _04918_ net263 _03325_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__and3_1
X_15735_ net1294 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12947_ net249 net2364 net321 vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XANTENNA__14529__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15666_ net1175 vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__inv_2
X_12878_ _07578_ net330 net388 net2159 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14617_ net1237 vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__inv_2
X_11829_ net2462 net526 net443 _07308_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__a22o_1
X_15597_ net1144 vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17336_ net1392 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14548_ net1192 vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__inv_2
XANTENNA__09711__S1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13963__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11974__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267_ net1327 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_0_141_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xclkload102 clknet_leaf_156_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload102/X sky130_fd_sc_hd__clkbuf_4
X_14479_ net1273 vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11240__X _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload113 clknet_leaf_163_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload113/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16218_ clknet_leaf_39_wb_clk_i _01887_ _00447_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload124 clknet_leaf_142_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload124/X sky130_fd_sc_hd__clkbuf_4
Xclkload135 clknet_leaf_64_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload135/Y sky130_fd_sc_hd__clkinv_4
Xclkload146 clknet_leaf_71_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload146/Y sky130_fd_sc_hd__inv_6
X_17198_ clknet_leaf_69_wb_clk_i _02810_ _01427_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload157 clknet_leaf_99_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload157/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_168_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload168 clknet_leaf_81_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload168/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_168_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16149_ clknet_leaf_33_wb_clk_i _01818_ _00378_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09792__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14125__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _04576_ _04581_ net725 vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_109_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07922_ net1098 net1076 vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__or2_1
Xhold19 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[31\]
+ vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13327__B team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08201__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09336__A1_N net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__mux2_1
XANTENNA__12658__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ net724 _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08405_ net727 _04015_ net712 vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__o21a_1
X_09385_ _04992_ _04993_ _04994_ _04995_ net793 net813 vssd1 vssd1 vccd1 vccd1 _04996_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout524_A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1266_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08336_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[26\] team_04_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12611__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11965__A2 _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07995__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08267_ net778 _03877_ net762 vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout312_X net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_148_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08198_ net644 _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__B net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14116__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10160_ _05672_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 _06000_ vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _04612_ vssd1
+ vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__and2b_1
XANTENNA__10641__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__clkbuf_2
Xfanout1028 _03539_ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1039 net1042 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09207__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11038__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ team_04_WB.ADDR_START_VAL_REG\[31\] _03240_ vssd1 vssd1 vccd1 vccd1 _03241_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12801_ net236 net2320 net322 vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__mux2_1
XANTENNA__11980__B _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13781_ _07751_ _07754_ _07824_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__and3_1
XANTENNA__10877__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ _06355_ _06470_ _06475_ _06479_ _06481_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a2111o_2
XFILLER_0_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14349__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15520_ net1153 vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__inv_2
X_12732_ _07457_ net329 net400 net2214 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
XANTENNA__12850__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_187_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15451_ net1136 vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12663_ net247 net2427 net475 vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ net1292 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11614_ net754 _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__nand2_1
XANTENNA__11405__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ net1223 vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12602__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ _07563_ net480 net412 net1962 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17121_ clknet_leaf_67_wb_clk_i _02756_ _01350_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14333_ _03364_ _03373_ _03492_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.pixel_data
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_137_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11545_ _06273_ _06578_ _06668_ _06884_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17052_ clknet_leaf_46_wb_clk_i _00018_ _01281_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14264_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] _03442_
+ net820 vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__o21ai_1
X_11476_ net574 _06963_ _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ clknet_leaf_52_wb_clk_i _01679_ _00232_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_10427_ _06004_ _06005_ _06002_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__o21a_1
X_13215_ net87 team_04_WB.MEM_SIZE_REG_REG\[26\] net982 vssd1 vssd1 vccd1 vccd1 _01688_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08034__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14195_ _03365_ _03360_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14107__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13146_ _07580_ net381 net297 net2316 vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12669__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ net254 net2216 net302 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_163_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ net622 _05881_ _05882_ _05885_ net281 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__a311o_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08337__B2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16905_ clknet_leaf_99_wb_clk_i _02574_ _01134_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\]
+ sky130_fd_sc_hd__dfrtp_1
X_12028_ net2380 net518 _07467_ net458 vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XANTENNA__11219__Y _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__Y _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16836_ clknet_leaf_173_wb_clk_i _02505_ _01065_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08956__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17339__1395 vssd1 vssd1 vccd1 vccd1 _17339__1395/HI net1395 sky130_fd_sc_hd__conb_1
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09641__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ clknet_leaf_156_wb_clk_i _02436_ _00996_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13094__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17252__1312 vssd1 vssd1 vccd1 vccd1 _17252__1312/HI net1312 sky130_fd_sc_hd__conb_1
XFILLER_0_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13979_ _04471_ net266 net599 _03323_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__a31o_1
X_15718_ net1295 vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__inv_2
XANTENNA__12841__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16698_ clknet_leaf_37_wb_clk_i _02367_ _00927_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\]
+ sky130_fd_sc_hd__dfrtp_1
X_15795__14 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__inv_2
XFILLER_0_76_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15649_ net1177 vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13397__A1 team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09787__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09170_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[7\] net1010
+ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08499__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08121_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\]
+ net851 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux2_1
X_17319_ net1375 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12066__X _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11411__A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09088__A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08052_ _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12941__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__A3 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10383__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A3 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13537__A1_N net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_1
XANTENNA__09027__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ net1087 vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08885_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__mux2_1
XANTENNA__13872__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10686__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13085__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10697__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _04001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\]
+ net879 vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12832__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout906_A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_679 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11799__Y _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09368_ _04755_ net366 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13520__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09299_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11330_ team_04_WB.MEM_SIZE_REG_REG\[23\] _06513_ team_04_WB.MEM_SIZE_REG_REG\[24\]
+ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11321__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout896_X net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11261_ _06272_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_132_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12899__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10212_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__nand2_1
X_13000_ _07649_ net468 net310 net2073 vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ net706 _06660_ _06679_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__or3_2
X_10143_ _05704_ _05753_ _05705_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__a21boi_1
XANTENNA__12115__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10074_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__inv_2
XANTENNA_input35_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ net1139 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13902_ _03274_ _03277_ net2569 net1066 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11991__A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14882_ net1265 vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__inv_2
X_16621_ clknet_leaf_28_wb_clk_i _02290_ _00850_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\]
+ sky130_fd_sc_hd__dfrtp_1
X_13833_ _02899_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__or2_1
XANTENNA__13076__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16552_ clknet_leaf_160_wb_clk_i _02221_ _00781_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11626__A1 _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ net1002 _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__or2_1
X_10976_ _04474_ _06464_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15503_ net1195 vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12715_ net1912 net407 net347 _07397_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16483_ clknet_leaf_122_wb_clk_i _02152_ _00712_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\]
+ sky130_fd_sc_hd__dfrtp_1
X_13695_ _03057_ _03084_ _03054_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15434_ net1106 vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12646_ _07617_ net490 net410 net1775 vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09400__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11502__Y _06991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10546__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ net1110 vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12577_ _07544_ net482 net416 net1759 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a22o_1
XANTENNA__12327__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ clknet_leaf_106_wb_clk_i _02739_ _01333_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14316_ net1087 _03472_ _03475_ net1089 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__o211ai_1
Xwire250 _07396_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_152_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _05460_ _06401_ _06884_ _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_113_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15296_ net1210 vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\] vssd1 vssd1
+ vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\] vssd1 vssd1
+ vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ clknet_leaf_17_wb_clk_i _02704_ _01264_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
X_14247_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] _03432_ vssd1
+ vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and2_1
XANTENNA__13000__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14542__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ net466 _06885_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__nor2_2
XFILLER_0_22_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12354__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ _03514_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ _07563_ net367 net294 net2071 vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__a22o_1
Xhold1008 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\] vssd1 vssd1
+ vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\] vssd1 vssd1
+ vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08670_ net720 _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__or2_1
XANTENNA__10668__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16819_ clknet_leaf_181_wb_clk_i _02488_ _01048_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12814__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__A1 _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09222_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12042__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout222_A _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08104_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__mux2_1
XANTENNA__12593__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ _04677_ _04683_ _04694_ net717 vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__a22o_2
XFILLER_0_142_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08035_ _03640_ net702 _03644_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__o21ai_2
Xinput80 wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold820 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\] vssd1 vssd1
+ vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12671__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput91 wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1131_A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold831 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\] vssd1 vssd1
+ vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\] vssd1 vssd1
+ vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\] vssd1 vssd1
+ vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold864 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\] vssd1 vssd1
+ vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\] vssd1 vssd1
+ vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout689_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold886 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\] vssd1 vssd1
+ vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[973\] vssd1 vssd1
+ vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ _05595_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__or2_1
XANTENNA__10108__A1 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
XANTENNA__13845__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout856_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11856__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08596__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__mux2_1
X_08799_ _04404_ _04409_ net723 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10830_ net643 _06316_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__and2_1
XANTENNA__12805__A0 _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ _05446_ _05469_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__nor2_2
XANTENNA__12281__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _07497_ net484 net425 net2235 vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08047__D net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13480_ net989 _02870_ _02867_ net994 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_62_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _04782_ net822 vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_62_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14022__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13230__A0 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08237__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ net2339 net434 _07636_ net523 vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10593__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08788__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08332__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__A3 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15150_ net1203 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__inv_2
XANTENNA__12584__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net214 net2514 net497 vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__mux2_1
X_17338__1394 vssd1 vssd1 vccd1 vccd1 _17338__1394/HI net1394 sky130_fd_sc_hd__conb_1
X_14101_ team_04_WB.EN_VAL_REG _06146_ _06153_ _03355_ vssd1 vssd1 vccd1 vccd1 net179
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_130_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08883__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ net593 net592 net638 net639 net543 net536 vssd1 vssd1 vccd1 vccd1 _06802_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15081_ net1132 vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__inv_2
X_12293_ _04783_ _05279_ _05406_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__or3_1
XANTENNA__14362__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17251__1311 vssd1 vssd1 vccd1 vccd1 _17251__1311/HI net1311 sky130_fd_sc_hd__conb_1
XFILLER_0_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12336__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14032_ net26 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1
+ vccd1 vccd1 _01554_ sky130_fd_sc_hd__o22a_1
X_11244_ _06454_ _06466_ _06472_ _06462_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__a211o_1
XANTENNA__09201__A2 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ net640 net595 net593 net592 net543 net536 vssd1 vssd1 vccd1 vccd1 _06664_
+ sky130_fd_sc_hd__mux4_1
X_10126_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] _05405_ _05407_
+ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or3_1
XANTENNA__08960__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15983_ clknet_leaf_51_wb_clk_i _01659_ _00212_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10057_ _03494_ _03783_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
X_14934_ net1228 vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13049__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14865_ net1265 vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload0_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16604_ clknet_leaf_126_wb_clk_i _02273_ _00833_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\]
+ sky130_fd_sc_hd__dfrtp_1
X_13816_ net992 _03203_ _03206_ net989 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_158_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14796_ net1121 vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16535_ clknet_leaf_167_wb_clk_i _02204_ _00764_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\]
+ sky130_fd_sc_hd__dfrtp_1
X_13747_ net999 _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ _06437_ _06446_ _06447_ _06431_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__a22o_1
XANTENNA__14537__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16466_ clknet_leaf_9_wb_clk_i _02135_ _00695_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13678_ _07116_ net274 _07693_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10784__B _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09130__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13221__A0 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15417_ net1251 vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12629_ _07600_ net485 net409 net1719 vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
X_16397_ clknet_leaf_40_wb_clk_i _02066_ _00626_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[370\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12024__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_171_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_171_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12575__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13772__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15348_ net1227 vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__inv_2
XANTENNA__11783__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[6\]
+ vssd1 vssd1 vccd1 vccd1 net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold116 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[11\]
+ vssd1 vssd1 vccd1 vccd1 net1553 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ net1196 vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__inv_2
Xhold127 net159 vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[22\] vssd1
+ vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\] vssd1 vssd1
+ vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ clknet_leaf_38_wb_clk_i _02687_ _01247_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09366__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09840_ _04669_ _05443_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__nor2_1
Xfanout607 net609 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
Xfanout618 net619 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10305__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout629 _04892_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12223__C net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09771_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\]
+ net962 vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08722_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XANTENNA__11838__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13335__B team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11136__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12263__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12666__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_A _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout437_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08562__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10813__A2 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09040__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09205_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13763__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__mux2_1
XANTENNA__13763__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11774__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09067_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12318__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ _03597_ _03616_ _03619_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__and3_1
Xhold650 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\] vssd1 vssd1
+ vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__B2 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09814__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\] vssd1 vssd1
+ vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold672 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\] vssd1 vssd1
+ vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\] vssd1 vssd1
+ vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold694 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\] vssd1 vssd1
+ vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13279__A0 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _04556_ _04559_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ net611 _07397_ net474 net316 net2164 vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_86_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ net655 net249 vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__and2_1
XANTENNA__10501__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14650_ net1146 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__inv_2
X_11862_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net270 net267 vssd1 vssd1 vccd1
+ vccd1 _07337_ sky130_fd_sc_hd__a21o_1
XFILLER_0_170_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ _02982_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__or2_1
XFILLER_0_169_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10813_ _04193_ net658 _06282_ _06300_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ net1178 vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08458__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14357__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11793_ net652 net217 vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08553__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16320_ clknet_leaf_136_wb_clk_i _01989_ _00549_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ _06858_ net272 net709 vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10744_ _06232_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16251_ clknet_leaf_101_wb_clk_i _01920_ _00480_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\]
+ sky130_fd_sc_hd__dfrtp_1
X_13463_ _03509_ _02852_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ net1626 net1017 net1013 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1
+ vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08305__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ net1218 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12557__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12414_ net521 net603 _07334_ net433 net1608 vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16182_ clknet_leaf_17_wb_clk_i _01851_ _00411_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\]
+ sky130_fd_sc_hd__dfrtp_1
X_13394_ _07766_ _07819_ _07818_ _07816_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15188__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ net1147 vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__inv_2
X_12345_ net233 net670 vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07984__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15064_ net1222 vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__inv_2
X_12276_ net261 net674 vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14015_ net1440 net1069 _03343_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__a21o_1
X_11227_ _06714_ _06715_ net557 vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__mux2_1
XANTENNA__10125__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14820__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08933__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__A net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_156_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_156_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11158_ net557 _05474_ _06642_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_147_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__A1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_147_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ _05718_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__nand2b_1
X_15966_ clknet_leaf_59_wb_clk_i _01642_ _00195_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_11089_ _06571_ _06577_ net562 vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__mux2_1
XANTENNA__09125__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14917_ net1109 vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire238_A _07313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ clknet_leaf_99_wb_clk_i _01574_ _00124_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_159_Right_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14848_ net1213 vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12339__X _07614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12245__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ net1126 vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__inv_2
XANTENNA__10795__A _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_173_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16518_ clknet_leaf_17_wb_clk_i _02187_ _00747_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[491\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16449_ clknet_leaf_141_wb_clk_i _02118_ _00678_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__S net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11756__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12234__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout404 _07664_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__buf_6
Xfanout415 _07660_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__buf_6
Xfanout426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_8
Xfanout437 net444 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12720__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _03634_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__o21ai_2
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__clkbuf_4
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_2
XANTENNA__12521__Y _07658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_A _07674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12250__A _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09035__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08705_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__mux2_1
X_09685_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__mux2_1
XANTENNA__13681__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1296_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_169_Left_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17337__1393 vssd1 vssd1 vccd1 vccd1 _17337__1393/HI net1393 sky130_fd_sc_hd__conb_1
X_08636_ net639 _04245_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__or2_1
XANTENNA__08874__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17250__1310 vssd1 vssd1 vccd1 vccd1 _17250__1310/HI net1310 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_81_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12787__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08498_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _06034_ _06035_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__mux2_1
X_10391_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__inv_2
XANTENNA__10644__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1__f_wb_clk_i_X clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12130_ net219 net2435 net511 vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12061_ net1975 net353 _07485_ net448 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\] vssd1 vssd1
+ vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold491 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\] vssd1 vssd1
+ vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ team_04_WB.MEM_SIZE_REG_REG\[5\] _06500_ vssd1 vssd1 vccd1 vccd1 _06501_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_25_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12711__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08915__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16236__CLK clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15820_ clknet_leaf_89_wb_clk_i _01497_ _00047_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_4
Xfanout971 net972 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_2
Xfanout982 net983 vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_4
Xfanout993 _07690_ vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_2
XANTENNA__10599__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15751_ net1269 vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__inv_2
X_12963_ net601 _07290_ net468 net314 net1681 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a32o_1
XANTENNA__11278__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13672__B1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1180 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\] vssd1 vssd1
+ vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14702_ net1198 vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__inv_2
Xhold1191 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\] vssd1 vssd1
+ vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07382_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15682_ net1256 vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__inv_2
X_12894_ _07596_ net333 net384 net1824 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ net1132 vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11845_ net758 _05871_ net697 _04331_ net693 vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__a221o_1
XANTENNA_output104_A net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13975__A1 _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12778__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14564_ net1176 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__inv_2
X_11776_ net705 _05790_ net690 _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__o211a_1
XANTENNA__08085__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11986__B1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16303_ clknet_leaf_186_wb_clk_i _01972_ _00532_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12319__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ net994 _02903_ _02905_ net989 vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o2bb2a_1
X_17283_ net1339 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10727_ _06214_ _06215_ net541 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__mux2_1
X_14495_ net1239 vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__inv_2
XANTENNA__11450__A2 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ clknet_leaf_164_wb_clk_i _01903_ _00463_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\]
+ sky130_fd_sc_hd__dfrtp_1
X_13446_ net1082 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 _07872_
+ sky130_fd_sc_hd__and2_1
X_10658_ net1525 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1
+ vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
Xclkload14 clknet_leaf_188_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_4
Xclkload25 clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/X sky130_fd_sc_hd__clkbuf_4
Xclkload36 clknet_leaf_181_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload36/X sky130_fd_sc_hd__clkbuf_4
X_16165_ clknet_leaf_5_wb_clk_i _01834_ _00394_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\]
+ sky130_fd_sc_hd__dfrtp_1
X_13377_ _07778_ _07780_ _07802_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__o21ba_1
Xclkload47 clknet_leaf_169_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload47/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ _06131_ net1534 net1023 vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__mux2_1
XANTENNA__12335__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload58 clknet_leaf_35_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload58/X sky130_fd_sc_hd__clkbuf_8
Xclkload69 clknet_leaf_50_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload69/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10781__C _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15116_ net1119 vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__inv_2
X_12328_ net2250 net501 _07608_ net451 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__a22o_1
X_16096_ clknet_leaf_140_wb_clk_i _01765_ _00325_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_149_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15047_ net1134 vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__inv_2
X_12259_ net2248 net504 _07572_ net446 vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_166_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12702__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12070__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16998_ clknet_leaf_20_wb_clk_i _02667_ _01227_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12466__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ clknet_leaf_43_wb_clk_i _01626_ _00176_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08765__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _05077_ _05078_ _05079_ _05080_ net835 net745 vssd1 vssd1 vccd1 vccd1 _05081_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08694__S net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08421_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__mux2_1
XANTENNA__12218__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12769__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08352_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\]
+ net862 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08283_ net752 _03893_ _03725_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a21o_2
XFILLER_0_116_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12944__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload8 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_8
XFILLER_0_15_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_138_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08282__X _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout302_A net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08070__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12154__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08869__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout212 _07258_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
Xfanout223 net225 vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_2
XANTENNA_fanout671_A _07589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net235 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout245 _07333_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_2
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09806_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_2
X_07998_ _03601_ _03603_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__and4_1
Xfanout289 _06526_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_2_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ _05344_ _05345_ _05346_ _05347_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_2_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout936_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12457__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09668_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] net974 _05278_ vssd1 vssd1 vccd1
+ vccd1 _05279_ sky130_fd_sc_hd__o21a_4
XANTENNA__15999__Q team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_177_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08619_ _04226_ _04227_ _04228_ _04229_ net823 net733 vssd1 vssd1 vccd1 vccd1 _04230_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10639__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\]
+ net957 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08508__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _06500_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__or2_1
XFILLER_0_166_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08109__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11968__B1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__A2 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _05336_ net548 net361 vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ net1082 team_04_WB.MEM_SIZE_REG_REG\[28\] vssd1 vssd1 vccd1 vccd1 _07726_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10512_ team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] net1094 net1054 vssd1 vssd1 vccd1
+ vccd1 _06080_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14280_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] _03452_
+ net821 vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11492_ net576 _06702_ _06948_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_98_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ net70 team_04_WB.MEM_SIZE_REG_REG\[10\] net984 vssd1 vssd1 vccd1 vccd1 _01672_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13185__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _06020_
+ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12393__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input65_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _07598_ net369 net290 net1593 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__a22o_1
X_10374_ _05720_ _05744_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_55_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ net2416 net354 _07511_ net453 vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__a22o_1
X_13093_ _07525_ net377 net300 net1867 vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__a22o_1
XANTENNA__12145__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08779__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16921_ clknet_leaf_152_wb_clk_i _02590_ _01150_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\]
+ sky130_fd_sc_hd__dfrtp_1
X_12044_ net2428 net517 _07475_ net453 vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16852_ clknet_leaf_3_wb_clk_i _02521_ _01081_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13612__A2_N net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout790 net799 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_161_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16783_ clknet_leaf_190_wb_clk_i _02452_ _01012_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13995_ _04864_ net263 _03325_ _03332_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_161_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15734_ net1295 vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__inv_2
XANTENNA__12999__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ net252 net2575 net318 vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09403__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15665_ net1175 vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__inv_2
X_12877_ _07577_ net328 net389 net2135 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14616_ net1207 vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__inv_2
X_11828_ net651 net247 vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15596_ net1119 vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12049__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17335_ net1391 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547_ net1259 vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11759_ net700 _06190_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17266_ net1326 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14478_ net1159 vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload103 clknet_leaf_109_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_116_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ clknet_leaf_175_wb_clk_i _01886_ _00446_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[190\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload114 clknet_leaf_130_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__bufinv_16
X_13429_ net1082 team_04_WB.MEM_SIZE_REG_REG\[26\] vssd1 vssd1 vccd1 vccd1 _07855_
+ sky130_fd_sc_hd__nand2_1
Xclkload125 clknet_leaf_115_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__inv_8
X_17197_ clknet_leaf_80_wb_clk_i _02809_ _01426_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_2
Xclkload136 clknet_leaf_91_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload136/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_116_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12384__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__A1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload147 clknet_leaf_72_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload147/Y sky130_fd_sc_hd__inv_6
XANTENNA__11187__B2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload158 clknet_leaf_101_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload158/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload169 clknet_leaf_82_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload169/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_168_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ clknet_leaf_2_wb_clk_i _01817_ _00377_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_168_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_171_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_171_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_17336__1392 vssd1 vssd1 vccd1 vccd1 _17336__1392/HI net1392 sky130_fd_sc_hd__conb_1
XANTENNA__14125__A1 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13595__S net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16079_ clknet_leaf_186_wb_clk_i _01748_ _00308_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_08970_ _04577_ _04578_ _04579_ _04580_ net831 net747 vssd1 vssd1 vccd1 vccd1 _04581_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08689__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12136__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ _03527_ _03530_ _03533_ _03534_ net1077 vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__a221o_2
XFILLER_0_20_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11895__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08760__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput1 ACK_I vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
XANTENNA__12939__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12439__B2 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[708\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__mux2_1
XANTENNA__09313__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _05060_ _05061_ _05062_ _05063_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05064_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08404_ _04011_ _04012_ _04013_ _04014_ net824 net733 vssd1 vssd1 vccd1 vccd1 _04015_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ net765 _03938_ _03944_ _03926_ _03932_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a32o_2
XANTENNA__11414__A2 _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12674__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08815__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1161_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout517_A _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1259_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08266_ _03873_ _03874_ _03875_ _03876_ net788 net804 vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__07995__C net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08197_ _03783_ _03807_ net662 vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__mux2_2
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12914__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14116__A1 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout886_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14116__B2 team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__Y _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12127__A0 _07246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08599__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10090_ _04612_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] vssd1
+ vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nand2b_1
Xfanout1007 _03653_ vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_2
Xfanout1018 _06176_ vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_2
Xfanout1029 _03539_ vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09543__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ net247 net2392 net322 vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13780_ net707 _06781_ net273 _07697_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__o31ai_1
X_10992_ net593 _06339_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09223__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ _07456_ net327 net400 net2052 vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15450_ net1142 vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ net240 net2522 net476 vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08915__X _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14401_ net1289 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11613_ _06204_ _07091_ _07095_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__o22a_2
XFILLER_0_136_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15381_ net1215 vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__inv_2
XANTENNA__10893__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _07562_ net483 net413 net2194 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__a22o_1
X_17120_ clknet_leaf_67_wb_clk_i _02755_ _01349_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14332_ _03485_ _03491_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08282__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11544_ net626 _05084_ net358 _07032_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17051_ clknet_leaf_46_wb_clk_i _00007_ _01280_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13158__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] _03442_
+ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ net568 _06803_ _06251_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12366__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ clknet_leaf_50_wb_clk_i _01678_ _00231_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_13214_ net88 team_04_WB.MEM_SIZE_REG_REG\[27\] net983 vssd1 vssd1 vccd1 vccd1 _01689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10426_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] _06001_
+ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__nand2_1
XANTENNA__08034__A1 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12905__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194_ net2651 _03371_ _03402_ _03534_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11220__C _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13145_ _07579_ net372 net294 net1922 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10357_ _05748_ _05945_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_111_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10392__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ net243 net2414 net302 vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__mux2_1
XANTENNA__08302__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13866__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ net622 _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__nor2_1
X_16904_ clknet_leaf_116_wb_clk_i _02573_ _01133_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\]
+ sky130_fd_sc_hd__dfrtp_1
X_12027_ net257 net684 vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__and2_1
XFILLER_0_174_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ clknet_leaf_124_wb_clk_i _02504_ _01064_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13618__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ clknet_leaf_142_wb_clk_i _02435_ _00995_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13978_ net144 net1070 vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09133__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15717_ net1295 vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__inv_2
X_12929_ net226 net2323 net318 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10301__C1 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16697_ clknet_leaf_152_wb_clk_i _02366_ _00926_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_124_Left_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15648_ net1180 vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15579_ net1114 vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08120_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\]
+ net851 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__mux2_1
X_17318_ net1374 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13149__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__nand2_4
X_17249_ net1309 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10368__C1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _04560_ _04561_ _04562_ _04563_ net837 net748 vssd1 vssd1 vccd1 vccd1 _04564_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12242__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ net1088 vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11868__C1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__mux2_1
XANTENNA__12669__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__X _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14282__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\]
+ net879 vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_861 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout801_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09367_ _04921_ _04922_ _04977_ _04867_ _04814_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_118_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_X net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12596__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08318_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[90\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__mux2_1
X_09298_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08249_ _03842_ _03848_ _03859_ net718 vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__a22o_4
XFILLER_0_160_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ net555 _06247_ _06571_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_132_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08470__X _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _03496_ net1055 _05816_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09764__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _06660_ _06679_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__nor2_1
XANTENNA__09218__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ _05707_ _05709_ _05751_ _05706_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput190 net190 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__buf_2
XANTENNA__15744__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _04274_ vssd1
+ vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or2_1
X_14950_ net1103 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__inv_2
X_13901_ _03148_ _03192_ _03243_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a21o_1
XANTENNA_input28_A DAT_I[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ net1188 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__inv_2
XANTENNA__10888__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ _03210_ _03219_ _03209_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a21o_1
X_16620_ clknet_leaf_112_wb_clk_i _02289_ _00849_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\]
+ sky130_fd_sc_hd__dfrtp_1
X_16551_ clknet_leaf_21_wb_clk_i _02220_ _00780_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13763_ net992 _03151_ _03153_ net989 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ _04528_ _06291_ net658 vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17335__1391 vssd1 vssd1 vccd1 vccd1 _17335__1391/HI net1391 sky130_fd_sc_hd__conb_1
XFILLER_0_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15502_ net1203 vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__inv_2
X_12714_ net2264 net404 net330 _07391_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16482_ clknet_leaf_146_wb_clk_i _02151_ _00711_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14025__B1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ _03057_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_167_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08792__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15433_ net1135 vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__inv_2
XANTENNA__09127__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12645_ _07616_ net487 net410 net1602 vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ net1187 vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__inv_2
X_12576_ _07543_ net480 net416 net1682 vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12327__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ net1088 _03473_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21o_1
X_17103_ clknet_leaf_106_wb_clk_i _02738_ _01332_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11527_ net566 _06872_ _06533_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_29_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15295_ net1249 vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire284 _06756_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_1
X_17034_ clknet_leaf_162_wb_clk_i _02703_ _01263_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
X_14246_ _03432_ net819 _03431_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__and3b_1
Xhold309 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] vssd1 vssd1
+ vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11458_ net566 _06741_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nor2_1
XANTENNA__08821__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1058 _05991_
+ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a21bo_1
X_14177_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _03389_
+ _03392_ _03378_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[4\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10562__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11389_ net287 _06874_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__and3_1
XANTENNA__12343__A _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13128_ _07562_ net374 net295 net2322 vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_12__f_wb_clk_i clknet_3_6_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12062__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ net215 net2413 net304 vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__mux2_1
Xhold1009 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\] vssd1 vssd1
+ vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12511__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16818_ clknet_leaf_8_wb_clk_i _02487_ _01047_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_132_Left_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16749_ clknet_leaf_29_wb_clk_i _02418_ _00978_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09798__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07900__A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09221_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12578__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__mux2_1
XANTENNA__12042__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08207__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08103_ _03710_ _03711_ _03712_ _03713_ net791 net812 vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12952__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _04688_ _04693_ net728 vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout215_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_141_Left_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08034_ _03640_ net702 _03644_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o21a_1
Xinput70 wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput81 wbs_dat_i[20] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold810 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\] vssd1 vssd1
+ vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\] vssd1 vssd1
+ vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 wbs_dat_i[30] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_1
Xhold832 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\] vssd1 vssd1
+ vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\] vssd1 vssd1
+ vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\] vssd1 vssd1
+ vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\] vssd1 vssd1
+ vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\] vssd1 vssd1
+ vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold887 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\] vssd1 vssd1
+ vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_71 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold898 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\] vssd1 vssd1
+ vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ net589 _05005_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08936_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
XANTENNA__10108__A2 _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08867_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_150_Left_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout849_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08178__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08798_ _04405_ _04406_ _04407_ _04408_ net829 net743 vssd1 vssd1 vccd1 vccd1 _04409_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_28_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11316__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10760_ _05446_ _05464_ _05470_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__or3_1
XANTENNA__12281__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ _05005_ _05029_ net665 vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__mux2_2
XFILLER_0_164_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10691_ net1605 net711 _06180_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
XANTENNA__12428__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12569__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12430_ net653 net607 net231 vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__and3_1
XFILLER_0_164_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08237__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10044__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ net212 net2461 net497 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__mux2_1
XANTENNA__08332__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14643__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ team_04_WB.MEM_SIZE_REG_REG\[0\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[0\]
+ net1004 vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__o221a_1
XANTENNA__11792__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _03891_ net642 net640 net595 net543 net535 vssd1 vssd1 vccd1 vccd1 _06801_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15080_ net1118 vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__inv_2
X_12292_ net822 _04782_ _05280_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__and3b_4
X_14031_ team_04_WB.instance_to_wrap.BUSY_O net1063 team_04_WB.instance_to_wrap.wb_manage.prev_BUSY_O
+ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__or3b_1
X_11243_ net753 _06729_ _06731_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12163__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ net535 _06661_ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10125_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _05342_ vssd1
+ vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15982_ clknet_leaf_47_wb_clk_i _01658_ _00211_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_10056_ _03494_ _03783_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor2_1
X_14933_ net1201 vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__inv_2
XANTENNA__10411__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ net1165 vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ clknet_leaf_100_wb_clk_i _02272_ _00832_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\]
+ sky130_fd_sc_hd__dfrtp_1
X_13815_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] _05824_ net1099
+ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14795_ net1162 vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14818__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_158_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13746_ _07692_ _03136_ _03134_ net995 vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16534_ clknet_leaf_11_wb_clk_i _02203_ _00763_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\]
+ sky130_fd_sc_hd__dfrtp_1
X_10958_ net632 _06430_ _06434_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11480__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ team_04_WB.ADDR_START_VAL_REG\[2\] _03066_ vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__xor2_1
X_16465_ clknet_leaf_181_wb_clk_i _02134_ _00694_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ _06376_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09899__C_N _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ _07599_ net481 net408 net1699 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a22o_1
X_15416_ net1205 vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12024__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16396_ clknet_leaf_120_wb_clk_i _02065_ _00625_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_171_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15347_ net1232 vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_171_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13772__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _07526_ net485 net417 net1828 vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22o_1
XANTENNA__14553__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11783__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09647__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12980__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15278_ net1198 vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__inv_2
Xhold106 net156 vssd1 vssd1 vccd1 vccd1 net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\] vssd1 vssd1
+ vccd1 vccd1 net1554 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[25\] vssd1
+ vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03422_ sky130_fd_sc_hd__and3_1
Xhold139 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[14\]
+ vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ clknet_leaf_178_wb_clk_i _02686_ _01246_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_644 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12732__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 net609 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__buf_2
Xfanout619 _05660_ vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08721_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__mux2_1
Xfanout1190 net1193 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11417__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__mux2_1
XANTENNA__09227__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11136__B _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ net592 _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12947__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_152_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12263__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08726__A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09321__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08562__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12248__A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout332_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1074_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__mux2_1
XANTENNA__08314__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12682__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11774__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11774__B2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09066_ net723 _04676_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08017_ _03615_ _03622_ net754 vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__or3_2
Xhold640 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\] vssd1 vssd1
+ vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\] vssd1 vssd1
+ vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 net108 vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12723__B1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17334__1390 vssd1 vssd1 vccd1 vccd1 _17334__1390/HI net1390 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_38_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\] vssd1 vssd1
+ vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\] vssd1 vssd1
+ vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold695 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\] vssd1 vssd1
+ vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09968_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__inv_2
X_08919_ net636 _04528_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09578__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08400__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ _03697_ _03753_ _03721_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or3b_1
XANTENNA__11829__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12430__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net695 _07008_ _07395_ net616 vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__a211oi_2
XANTENNA__11327__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ net758 _05888_ net697 _04441_ net694 vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a221o_1
XANTENNA__14323__S0 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_X net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13600_ team_04_WB.ADDR_START_VAL_REG\[12\] _02989_ vssd1 vssd1 vccd1 vccd1 _02991_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_64_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _06282_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14580_ net1192 vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08458__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ net693 _06651_ _07276_ net615 vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_0_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _02910_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08553__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10743_ _06230_ _06231_ net537 vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11062__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16250_ clknet_leaf_40_wb_clk_i _01919_ _00479_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\]
+ sky130_fd_sc_hd__dfrtp_1
X_13462_ _03509_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__or2_1
XANTENNA_input95_A wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ net1504 net1018 net1014 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1
+ vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15201_ net1169 vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__inv_2
XANTENNA__11997__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12413_ net522 net604 _07328_ net433 net1610 vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a32o_1
XANTENNA__08305__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16181_ clknet_leaf_33_wb_clk_i _01850_ _00410_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\]
+ sky130_fd_sc_hd__dfrtp_1
X_13393_ _07764_ _07818_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__nand2_1
XANTENNA__11765__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15132_ net1148 vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__inv_2
XANTENNA__12962__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12344_ net2245 net501 _07616_ net452 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ net1231 vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__inv_2
XANTENNA__07984__A3 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08069__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12275_ net2541 net506 _07580_ net458 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a22o_1
XANTENNA__12714__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ _05432_ net264 _03335_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__and3_1
X_11226_ net592 net639 net638 _04328_ net535 net545 vssd1 vssd1 vccd1 vccd1 _06715_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12190__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__B net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ _03892_ _03919_ _06257_ _06645_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _03724_ _03893_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__a21o_1
XANTENNA__17192__Q team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15965_ clknet_leaf_69_wb_clk_i _01641_ _00194_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11088_ _06576_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__inv_2
XANTENNA__11237__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _05557_ _05649_ _05558_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__o21ai_1
X_14916_ net1189 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15896_ clknet_leaf_99_wb_clk_i _01573_ _00123_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_72_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14847_ net1248 vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_19_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12245__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778_ net1147 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_173_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16517_ clknet_leaf_5_wb_clk_i _02186_ _00746_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_173_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13729_ team_04_WB.ADDR_START_VAL_REG\[10\] _03117_ vssd1 vssd1 vccd1 vccd1 _03120_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__13993__A2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_128_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16448_ clknet_leaf_139_wb_clk_i _02117_ _00677_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16379_ clknet_leaf_104_wb_clk_i _02048_ _00608_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12355__X _07622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11756__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout405 _07664_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_4
Xfanout416 net419 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_8
X_09822_ net666 _05408_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__or2_1
Xfanout427 _07656_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_4
XANTENNA__12090__X _07500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__X _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 net444 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
Xfanout449 _07252_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09316__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__mux2_1
XANTENNA__08220__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ net773 _04308_ _04314_ net762 vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o211a_1
XANTENNA__13130__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ net730 _05288_ net715 vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08688__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08635_ _04245_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__inv_2
XANTENNA__11692__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_167_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_96_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12677__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11434__X _06923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1289_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09051__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[759\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout714_A net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08860__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13197__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12944__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10390_ _05527_ _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09049_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12060_ net211 net677 vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__and2_1
Xhold470 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\] vssd1 vssd1
+ vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold481 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\] vssd1 vssd1
+ vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout969_X net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ team_04_WB.MEM_SIZE_REG_REG\[4\] team_04_WB.MEM_SIZE_REG_REG\[3\] team_04_WB.MEM_SIZE_REG_REG\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and3_1
Xhold492 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\] vssd1 vssd1
+ vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09226__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 net972 vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
Xfanout961 net962 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_2
XANTENNA__08130__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout972 _03555_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__clkbuf_2
Xfanout983 net985 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__clkbuf_4
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_2
XANTENNA__10599__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13121__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ net1277 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__inv_2
X_12962_ net603 _07284_ net470 net315 net1611 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__a32o_1
XANTENNA__12475__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11278__A3 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[849\] vssd1 vssd1
+ vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A DAT_I[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10486__A1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ net1210 vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__inv_2
X_11913_ net2098 net526 net439 _07381_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a22o_1
Xhold1181 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\] vssd1 vssd1
+ vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1192 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\] vssd1 vssd1
+ vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15681_ net1281 vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__inv_2
X_12893_ _07595_ net341 net386 net1808 vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ net2230 net526 net436 _07321_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
X_14632_ net1117 vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__inv_2
XANTENNA__08366__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12159__Y _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14563_ net1176 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09723__S0 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ net687 _07260_ _07261_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13975__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11986__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ clknet_leaf_26_wb_clk_i _01971_ _00531_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\]
+ sky130_fd_sc_hd__dfrtp_1
X_13514_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _05837_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__mux2_1
X_10726_ net589 net626 net551 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__mux2_1
X_17282_ net1338 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XANTENNA_input98_X net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14494_ net1251 vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11450__A3 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13188__B1 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ net1083 team_04_WB.MEM_SIZE_REG_REG\[29\] vssd1 vssd1 vccd1 vccd1 _07871_
+ sky130_fd_sc_hd__nor2_1
X_16233_ clknet_leaf_121_wb_clk_i _01902_ _00462_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\]
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ net1524 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1
+ vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a22o_1
XANTENNA__11520__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload15 clknet_leaf_189_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload26 clknet_leaf_170_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__bufinv_16
X_13376_ _07783_ _07801_ _07781_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__o21a_1
Xclkload37 clknet_leaf_183_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ clknet_leaf_21_wb_clk_i _01833_ _00393_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\]
+ sky130_fd_sc_hd__dfrtp_1
X_10588_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[4\]
+ _06130_ net1050 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12335__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload48 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload48/X sky130_fd_sc_hd__clkbuf_8
Xclkload59 clknet_leaf_36_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
X_12327_ net258 net671 vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15115_ net1160 vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16095_ clknet_leaf_156_wb_clk_i _01764_ _00324_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_149_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15046_ net1105 vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__inv_2
X_12258_ _07349_ net673 vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__and2_1
X_11209_ _06614_ _06617_ net562 vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__mux2_1
XANTENNA__11519__X _07008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12189_ net244 net650 vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11910__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire250_A _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16997_ clknet_leaf_185_wb_clk_i _02666_ _01226_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12070__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15948_ clknet_leaf_46_wb_clk_i _01625_ _00175_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12466__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08765__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15879_ clknet_leaf_79_wb_clk_i _01556_ _00106_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__dfrtp_1
X_08420_ net640 _04029_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__xor2_1
XANTENNA__12218__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08351_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\]
+ net862 vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[27\] team_04_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__mux2_4
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload9 clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__13179__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_964 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_93_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12926__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08215__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14128__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10401__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09835__A _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout497_A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13357__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 _07258_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__buf_1
XFILLER_0_100_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout224 net225 vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_1
Xfanout246 _07320_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09805_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\]
+ net890 vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A DAT_I[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 _07241_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_31_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout279 _05524_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_4
X_07997_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout664_A net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09736_ _03508_ _03651_ net1007 _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a311o_1
XANTENNA__12457__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[9\] net1009
+ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout831_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1194_X net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout929_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08618_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
X_09598_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08549_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__mux2_1
XANTENNA__08508__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__A1 _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11968__B2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09181__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ net578 _07004_ _07047_ _07048_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__o22a_1
XANTENNA__11432__A3 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ _06079_ net1823 net1023 vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11491_ _06692_ _06887_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12436__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ net71 team_04_WB.MEM_SIZE_REG_REG\[11\] net984 vssd1 vssd1 vccd1 vccd1 _01673_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12917__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10442_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _06020_
+ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_98_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08125__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12393__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14119__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13590__B1 team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13161_ _07597_ net374 net291 net1917 vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__a22o_1
X_10373_ _05597_ _05598_ _05620_ net617 vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12112_ net224 net678 vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input58_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _07524_ net376 net300 net1943 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a22o_1
X_16920_ clknet_leaf_150_wb_clk_i _02589_ _01149_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\]
+ sky130_fd_sc_hd__dfrtp_1
X_12043_ net233 net683 vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12171__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12696__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16851_ clknet_leaf_183_wb_clk_i _02520_ _01080_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout791 net799 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_4_14__f_wb_clk_i_A clknet_3_7_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16782_ clknet_leaf_30_wb_clk_i _02451_ _01011_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_161_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ net137 net1065 vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_161_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ net1295 vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__inv_2
XANTENNA__11656__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ _07385_ net2429 net318 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
X_15664_ net1173 vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__inv_2
X_12876_ _07576_ net339 net389 net2149 vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14615_ net1223 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11827_ net689 _06680_ _07306_ net613 vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__o211a_2
X_15595_ net1159 vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17313__1369 vssd1 vssd1 vccd1 vccd1 _17313__1369/HI net1369 sky130_fd_sc_hd__conb_1
XFILLER_0_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ net1390 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_139_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14546_ net1259 vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12081__B1 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11758_ net652 net211 vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10709_ _06189_ _06196_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__or2_4
X_17265_ net1325 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XANTENNA__10565__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11689_ _04142_ _06248_ net362 _04141_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__a221o_1
X_14477_ net1159 vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12908__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload104 clknet_leaf_110_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload104/X sky130_fd_sc_hd__clkbuf_8
X_16216_ clknet_leaf_153_wb_clk_i _01885_ _00445_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\]
+ sky130_fd_sc_hd__dfrtp_1
X_13428_ _07737_ _07853_ _07734_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_116_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload115 clknet_leaf_132_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload115/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17196_ clknet_leaf_78_wb_clk_i _02808_ _01425_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkload126 clknet_leaf_116_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload126/X sky130_fd_sc_hd__clkbuf_8
Xclkload137 clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload137/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload148 clknet_leaf_73_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload148/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload159 clknet_leaf_102_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload159/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_168_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13359_ _07783_ _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__or2_1
X_16147_ clknet_leaf_182_wb_clk_i _01816_ _00376_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_168_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14125__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16078_ clknet_leaf_30_wb_clk_i _01747_ _00307_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07920_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\] team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__and2b_1
XANTENNA__09001__A1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15029_ net1211 vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__inv_2
XANTENNA__11895__B1 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15392__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 DAT_I[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12439__A2 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\]
+ net882 vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__mux2_1
XANTENNA__13734__A2_N net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08403_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__mux2_1
X_09383_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12955__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14061__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_136_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout245_A _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14736__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08334_ net765 _03938_ _03944_ _03926_ _03932_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08815__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12611__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08265_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\]
+ net930 vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07995__D net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12256__A _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08196_ net718 _03806_ _03795_ _03789_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14116__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1008 _03651_ vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_2
Xfanout1019 _06176_ vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09852__X _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11886__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_27_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09719_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[704\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__mux2_1
X_10991_ net593 _06339_ _06342_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ _07455_ net334 net401 net1906 vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XANTENNA__10310__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ net241 net2382 net475 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14052__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14400_ net1289 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _06718_ _06886_ _06948_ _06724_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12063__B1 _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15380_ net1236 vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__inv_2
X_12592_ _07561_ net485 net413 net2176 vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__a22o_1
XANTENNA__08644__A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14331_ _03519_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03486_ _03490_
+ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a41o_1
XFILLER_0_135_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11543_ _05086_ net365 net361 _05085_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_137_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14262_ _03442_ net820 _03441_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__and3b_1
X_17050_ clknet_leaf_38_wb_clk_i _02719_ _01279_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
X_11474_ net560 _06960_ _06961_ _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16001_ clknet_leaf_50_wb_clk_i _01677_ _00230_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[15\]
+ sky130_fd_sc_hd__dfrtp_4
X_13213_ net89 team_04_WB.MEM_SIZE_REG_REG\[28\] net983 vssd1 vssd1 vccd1 vccd1 _01690_
+ sky130_fd_sc_hd__mux2_1
X_10425_ _03514_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__and2_1
XANTENNA__09767__C1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ _03374_ _03375_ _03532_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_74_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14107__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ _07578_ net372 net294 net2628 vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__a22o_1
XANTENNA__09475__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ _05714_ _05716_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1111 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_11__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13075_ net255 net2296 net305 vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__mux2_1
X_10287_ _05757_ _05883_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13866__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ net2600 net517 _07466_ net442 vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
X_16903_ clknet_leaf_165_wb_clk_i _02572_ _01132_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11877__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13725__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16834_ clknet_leaf_147_wb_clk_i _02503_ _01063_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13618__A1 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16765_ clknet_leaf_131_wb_clk_i _02434_ _00994_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\]
+ sky130_fd_sc_hd__dfrtp_1
X_13977_ net1717 net1065 _03322_ net262 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a22o_1
XANTENNA__13094__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15716_ net1295 vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12928_ net227 net2374 net319 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__mux2_1
X_16696_ clknet_leaf_153_wb_clk_i _02365_ _00925_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12841__A2 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ net1180 vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__inv_2
X_12859_ _07559_ net340 net390 net2148 vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__a22o_1
XANTENNA__14043__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13460__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_791 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15578_ net1151 vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17317_ net1373 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14529_ net1193 vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__inv_2
XANTENNA__11801__B1 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ net1079 net1028 net1024 _03501_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__a31o_2
X_17248_ net1308 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_4_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap711 _06179_ vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__buf_4
X_17179_ clknet_leaf_92_wb_clk_i _02791_ _01408_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12109__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08952_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__mux2_1
X_07903_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\] vssd1 vssd1 vccd1 vccd1
+ _03518_ sky130_fd_sc_hd__inv_2
XANTENNA__11868__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ _04490_ _04491_ _04492_ _04493_ net788 net809 vssd1 vssd1 vccd1 vccd1 _04494_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11707__X _07196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09504_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[388\]
+ net880 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_wb_clk_i_X clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_116_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12832__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12685__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1271_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14034__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout627_A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ net627 _04973_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_23_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08317_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_40 net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_260 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08248_ _03853_ _03858_ net725 vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12348__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12899__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ net277 _05815_ _05813_ net1074 vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08403__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ _06673_ _06676_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _05709_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput180 net180 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput191 net191 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
XFILLER_0_101_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17312__1368 vssd1 vssd1 vccd1 vccd1 _17312__1368/HI net1368 sky130_fd_sc_hd__conb_1
X_10072_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] _04167_ vssd1
+ vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ net1689 net1066 _03275_ _03276_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a22o_1
X_14880_ net1213 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__inv_2
X_13831_ _03194_ _03199_ _03221_ _02948_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_159_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16550_ clknet_leaf_22_wb_clk_i _02219_ _00779_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\]
+ sky130_fd_sc_hd__dfrtp_1
X_13762_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] _05871_ net1100
+ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__mux2_1
X_10974_ _06459_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15501_ net1143 vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_139_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ net1863 net404 net328 _07386_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a22o_1
X_16481_ clknet_leaf_130_wb_clk_i _02150_ _00710_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ _03068_ _03082_ _03067_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_139_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_199 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15432_ net1117 vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__inv_2
XANTENNA__09127__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12644_ _07615_ net492 net411 net1802 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ _07542_ net485 net417 net2031 vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
X_15363_ net1168 vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11795__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17102_ clknet_leaf_104_wb_clk_i _02737_ _01331_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input80_X net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[21\]
+ _03357_ _03471_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[20\]
+ _03520_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ _06871_ _07014_ net576 vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__mux2_1
Xwire252 _07390_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_2
X_15294_ net1214 vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17033_ clknet_leaf_100_wb_clk_i _02702_ _01262_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
X_14245_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\]
+ _03428_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11457_ net566 _06742_ _06533_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__o21a_1
Xwire285 _07128_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__buf_1
XFILLER_0_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13000__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ net283 _05989_ _05990_ _05987_ net1058 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09409__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14176_ _03385_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08313__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _04586_ net364 _06272_ _06225_ _06876_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__o221a_1
XANTENNA__17195__Q team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10339_ net623 _05928_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nor2_1
X_13127_ _07561_ net369 net294 net2170 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__a22o_1
X_13058_ net213 net2563 net304 vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_X clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12009_ net239 net681 vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10798__B _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16817_ clknet_leaf_179_wb_clk_i _02486_ _01046_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\]
+ sky130_fd_sc_hd__dfrtp_1
X_16748_ clknet_leaf_110_wb_clk_i _02417_ _00977_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08983__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16679_ clknet_leaf_168_wb_clk_i _02348_ _00908_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08555__Y _04166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09220_ _04827_ _04828_ _04829_ _04830_ net786 net807 vssd1 vssd1 vccd1 vccd1 _04831_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08877__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08102_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09082_ _04689_ _04690_ _04691_ _04692_ net826 net742 vssd1 vssd1 vccd1 vccd1 _04693_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08033_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[31\] team_04_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__mux2_4
XFILLER_0_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput60 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
Xhold800 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\] vssd1 vssd1
+ vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10753__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput71 wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_4
Xhold811 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\] vssd1 vssd1
+ vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_1
XFILLER_0_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput93 wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__buf_1
Xhold822 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\] vssd1 vssd1
+ vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09319__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold833 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\] vssd1 vssd1
+ vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\] vssd1 vssd1
+ vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\] vssd1 vssd1
+ vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\] vssd1 vssd1
+ vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10210__C1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold877 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[512\] vssd1 vssd1
+ vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\] vssd1 vssd1
+ vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _05003_ _05005_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__nor2_1
Xhold899 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\] vssd1 vssd1
+ vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08935_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08866_ _04475_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__nand2_1
XANTENNA__09054__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout744_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08893__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ net718 _05028_ _05017_ _05016_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__o2bb2a_4
X_10690_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\] net711 _06180_
+ net2309 vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12428__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09349_ net731 _04953_ net715 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_134_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11777__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ net211 net2612 net496 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__mux2_1
XANTENNA__10044__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ net573 _06794_ _06799_ net581 vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__a211o_1
XANTENNA__11792__A2 _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12291_ net2545 net506 _07588_ net460 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12444__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14030_ team_04_WB.instance_to_wrap.BUSY_O team_04_WB.instance_to_wrap.wb_manage.prev_BUSY_O
+ net1061 vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__and3b_1
X_11242_ _06511_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__and2_1
XANTENNA__08133__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12163__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _06561_ _06563_ net535 vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07972__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input40_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _05405_ _05407_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__o21a_1
X_15981_ clknet_leaf_43_wb_clk_i _01657_ _00210_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10899__A net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _03836_ vssd1
+ vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__nand2_1
X_14932_ net1235 vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__inv_2
XANTENNA__11701__C1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14863_ net1199 vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__inv_2
XANTENNA__13049__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16602_ clknet_leaf_36_wb_clk_i _02271_ _00831_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\]
+ sky130_fd_sc_hd__dfrtp_1
X_13814_ net996 _03204_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__or2_1
X_14794_ net1106 vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16533_ clknet_leaf_35_wb_clk_i _02202_ _00762_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\]
+ sky130_fd_sc_hd__dfrtp_1
X_13745_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _05952_ net1102
+ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10957_ _06381_ _06441_ _06440_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13214__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10283__A2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ clknet_leaf_1_wb_clk_i _02133_ _00693_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11480__A1 _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ team_04_WB.ADDR_START_VAL_REG\[2\] _03066_ vssd1 vssd1 vccd1 vccd1 _03067_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_118_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08308__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10888_ _04723_ _06375_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415_ net1233 vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ _07598_ net479 net408 net2120 vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ clknet_leaf_23_wb_clk_i _02064_ _00624_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11810__X _07292_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12057__C _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15346_ net1244 vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08391__X _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08633__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12558_ _07525_ net482 net416 net1921 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_171_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12980__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _06533_ _06823_ _06887_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ net1199 vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__inv_2
Xhold107 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[27\]
+ vssd1 vssd1 vccd1 vccd1 net1544 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _07486_ net487 net426 net1669 vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold118 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[1\] vssd1
+ vssd1 vccd1 vccd1 net1555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 net122 vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17016_ clknet_leaf_150_wb_clk_i _02685_ _01245_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\]
+ sky130_fd_sc_hd__dfrtp_1
X_14228_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\] vssd1 vssd1 vccd1
+ vccd1 _03421_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14159_ _03371_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout609 net612 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XANTENNA__08978__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08720_ net769 net702 _04330_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12496__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1180 net1181 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__clkbuf_4
Xfanout1191 net1193 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_4
X_08651_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_157_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08582_ _04167_ _04192_ net663 vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__mux2_2
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09602__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10274__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08218__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12248__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09203_ net633 net590 vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__xor2_2
XFILLER_0_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311__1367 vssd1 vssd1 vccd1 vccd1 _17311__1367/HI net1367 sky130_fd_sc_hd__conb_1
XANTENNA_fanout325_A _07671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _04741_ _04742_ _04743_ _04744_ net832 net737 vssd1 vssd1 vccd1 vccd1 _04745_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12420__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12971__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ _04672_ _04673_ _04674_ _04675_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04676_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12264__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1234_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ _03618_ _03625_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__or2_1
Xhold630 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\] vssd1 vssd1
+ vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout694_A _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\] vssd1 vssd1
+ vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\] vssd1 vssd1
+ vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13920__B1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold663 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\] vssd1 vssd1
+ vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold674 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\] vssd1 vssd1
+ vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\] vssd1 vssd1
+ vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold696 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\] vssd1 vssd1
+ vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ _04557_ _04558_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout861_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ net636 _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__nand2_1
XANTENNA__10512__A team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09578__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09898_ net646 _03694_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__nand2_1
XANTENNA__12430__C net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ net705 _05884_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nor2_1
XANTENNA__14323__S1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _04245_ _06291_ _06298_ net658 vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ net704 _05803_ net689 _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_0_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout914_X net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ _02919_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__nor2_1
XANTENNA__10265__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _04328_ net591 net549 vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_101_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11462__B2 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13461_ _07697_ _07725_ _02849_ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a22o_1
X_10673_ net1540 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1
+ vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14654__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_173_Right_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15200_ net1211 vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__inv_2
XFILLER_0_164_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12412_ net519 net600 _07321_ net432 net1581 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a32o_1
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ clknet_leaf_6_wb_clk_i _01849_ _00409_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\]
+ sky130_fd_sc_hd__dfrtp_1
X_13392_ net1085 team_04_WB.MEM_SIZE_REG_REG\[12\] _07761_ _07817_ vssd1 vssd1 vccd1
+ vccd1 _07818_ sky130_fd_sc_hd__o22ai_1
XANTENNA_input88_A wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15131_ net1113 vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__inv_2
XANTENNA__12962__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ _07402_ net670 vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ net1228 vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__inv_2
X_12274_ net249 net675 vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_79_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08069__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10406__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14013_ net1532 net1069 _03342_ net264 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a22o_1
X_11225_ net642 net640 net595 net593 net544 net535 vssd1 vssd1 vccd1 vccd1 _06714_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10725__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12190__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ _03892_ _03919_ net362 vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o21a_1
XFILLER_0_101_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10107_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] _03724_ _03893_
+ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__and3_1
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15964_ clknet_leaf_69_wb_clk_i _01640_ _00193_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11087_ _06573_ _06575_ net541 vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__mux2_1
X_14915_ net1175 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__inv_2
X_10038_ net596 _04056_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_125_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09894__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15895_ clknet_leaf_35_wb_clk_i _01572_ _00122_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09894__B2 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14846_ net1217 vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__inv_2
XANTENNA__08827__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ net1235 vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12349__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ net2499 net529 net460 _07446_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16516_ clknet_leaf_168_wb_clk_i _02185_ _00745_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_173_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13728_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_173_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12650__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_165_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_165_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12068__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16447_ clknet_leaf_161_wb_clk_i _02116_ _00676_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[420\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13659_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] _03025_ vssd1
+ vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_140_Right_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12402__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16378_ clknet_leaf_38_wb_clk_i _02047_ _00607_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[351\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15329_ net1167 vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 _07664_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_6
Xfanout417 net419 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_4
X_09821_ _05414_ _05420_ _05431_ net719 vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__a22o_2
XANTENNA__09393__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 _07641_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_8
Xfanout439 net444 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12469__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ net778 _04313_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__or2_1
X_09683_ net724 _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__nor2_1
XANTENNA__10051__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__A2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ net661 _04243_ _04244_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__o21bai_4
XANTENNA__09332__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13969__B1 _03318_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08565_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1184_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08496_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__mux2_1
XANTENNA__12641__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13197__A1 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09117_ net702 _04725_ _04330_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1237_X net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__X _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09048_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold460 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\] vssd1 vssd1
+ vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold471 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\] vssd1 vssd1
+ vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net707 _06498_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__nor2_1
XANTENNA__11904__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold482 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\] vssd1 vssd1
+ vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold493 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\] vssd1 vssd1
+ vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08411__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__A0 net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_2
XANTENNA__13535__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__clkbuf_4
Xfanout962 net972 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_2
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_4
Xfanout984 net985 vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_4
Xfanout995 _07689_ vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _07629_ net470 net315 net1715 vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__a22o_1
XANTENNA__09876__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1160 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\] vssd1 vssd1
+ vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\] vssd1 vssd1
+ vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
X_14700_ net1121 vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__inv_2
Xhold1182 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\] vssd1 vssd1
+ vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ net656 _07380_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__and2_1
XANTENNA__10486__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ net1262 vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_142_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _07594_ net340 net386 net1674 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22o_1
XANTENNA__12880__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1193 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\] vssd1 vssd1
+ vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09242__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14631_ net1137 vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ net651 net246 vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11435__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562_ net1184 vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__inv_2
XANTENNA__12632__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ net758 _05793_ net697 _03836_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__a22o_1
XANTENNA__13975__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09723__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16301_ clknet_leaf_44_wb_clk_i _01970_ _00530_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13513_ net1092 _02903_ net1043 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11986__A2 _07057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17281_ net1337 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
X_10725_ net588 net580 net547 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__mux2_1
X_14493_ net1120 vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16232_ clknet_leaf_113_wb_clk_i _01901_ _00461_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\]
+ sky130_fd_sc_hd__dfrtp_1
X_13444_ _07859_ _07862_ _07865_ _07869_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ net1565 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1
+ vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11520__B _07008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload16 clknet_leaf_190_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__clkinvlp_4
X_16163_ clknet_leaf_116_wb_clk_i _01832_ _00392_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\]
+ sky130_fd_sc_hd__dfrtp_1
X_13375_ _07785_ _07800_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__nor2_1
X_10587_ team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] net1096 net1053 vssd1 vssd1 vccd1
+ vccd1 _06130_ sky130_fd_sc_hd__and3_1
Xclkload27 clknet_leaf_171_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload38 clknet_leaf_184_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload38/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_152_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload49 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__bufinv_16
X_15114_ net1105 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_77_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09765__X _05376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12326_ net2361 net500 _07607_ net446 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__a22o_1
X_16094_ clknet_leaf_142_wb_clk_i _01763_ _00323_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15045_ net1108 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12699__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ net2607 net506 _07571_ net459 vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XANTENNA__09417__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ net573 _06694_ _06696_ net585 vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__o211a_1
X_12188_ net2259 net508 _07535_ net447 vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12351__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_166_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11139_ _06625_ _06626_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__xnor2_1
X_16996_ clknet_leaf_169_wb_clk_i _02665_ _01225_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\]
+ sky130_fd_sc_hd__dfrtp_1
X_17310__1366 vssd1 vssd1 vccd1 vccd1 _17310__1366/HI net1366 sky130_fd_sc_hd__conb_1
XANTENNA__09941__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15947_ clknet_leaf_46_wb_clk_i _01624_ _00174_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09411__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__Y _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15878_ clknet_leaf_52_wb_clk_i _01555_ _00105_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12871__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14829_ net1210 vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ net728 _03954_ net713 vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o21a_1
XANTENNA__11426__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12623__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ _03872_ _03878_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__a22o_4
XFILLER_0_128_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10739__C_N _06226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09327__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 net216 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__buf_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout392_A _07672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11968__A1_N _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
Xfanout247 _07307_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_2
X_09804_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[193\]
+ net893 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout258 _07356_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_2
Xfanout269 net270 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
X_07996_ _03605_ _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_2_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ net1008 _03653_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\]
+ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_2_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09858__B2 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ net756 _03623_ _03636_ net740 vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12862__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09062__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08617_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout824_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _04155_ _04156_ _04157_ _04158_ net785 net801 vssd1 vssd1 vccd1 vccd1 _04159_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12614__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09086__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[30\]
+ _06078_ net1048 vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11490_ _06442_ _06977_ net465 vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__o21a_1
XFILLER_0_163_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08406__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire637 _04472_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12436__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10441_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06012_
+ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_98_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11276__S0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14932__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14119__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09794__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ _05528_ _05958_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__or2_1
X_13160_ _07596_ net369 net290 net1645 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ net2446 net354 _07510_ net454 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10__f_wb_clk_i clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_13091_ _07523_ net376 net300 net2012 vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ net2236 net517 _07474_ net453 vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XANTENNA__09237__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\] vssd1 vssd1
+ vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12171__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_144_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16850_ clknet_leaf_8_wb_clk_i _02519_ _01079_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_4
Xfanout792 net799 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
X_16781_ clknet_leaf_32_wb_clk_i _02450_ _01010_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\]
+ sky130_fd_sc_hd__dfrtp_1
X_13993_ net1449 net1064 _03331_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_161_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ net1293 vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__inv_2
XANTENNA__11656__A1 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ net254 net2595 net318 vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__mux2_1
XANTENNA__10700__A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08377__A net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15663_ net1173 vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__inv_2
X_12875_ _07575_ net345 net391 net2155 vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
XANTENNA_output207_A net207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14614_ net1221 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__inv_2
X_15810__29 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__inv_2
X_11826_ net686 _07305_ _07304_ _07303_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12605__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15594_ net1107 vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__inv_2
X_17333_ net1389 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14545_ net1260 vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11757_ net694 _06498_ _07245_ net615 vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__a211oi_4
XANTENNA__12081__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17264_ net1324 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
X_10708_ _06189_ _06196_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__nor2_4
XFILLER_0_154_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14476_ net1188 vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__inv_2
X_11688_ net594 _04139_ _06257_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__and3b_1
XANTENNA__12908__A1 _07610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16215_ clknet_leaf_161_wb_clk_i _01884_ _00444_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\]
+ sky130_fd_sc_hd__dfrtp_1
X_13427_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload105 clknet_leaf_111_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__bufinv_16
X_17195_ clknet_leaf_79_wb_clk_i _02807_ _01424_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10639_ net1515 team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__mux2_1
Xclkload116 clknet_leaf_134_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__13030__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload127 clknet_leaf_117_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__inv_8
Xclkload138 clknet_leaf_106_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload138/Y sky130_fd_sc_hd__inv_8
Xclkload149 clknet_leaf_76_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload149/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__09936__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16146_ clknet_leaf_7_wb_clk_i _01815_ _00375_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_13358_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] team_04_WB.MEM_SIZE_REG_REG\[5\]
+ _07778_ _07782_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_168_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ net242 net668 vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__and2_1
X_16077_ clknet_leaf_42_wb_clk_i _01746_ _00306_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _03517_ _07718_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15028_ net1214 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15673__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11895__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13097__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16979_ clknet_leaf_181_wb_clk_i _02648_ _01208_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput3 DAT_I[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_1
XANTENNA__13193__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__mux2_1
XANTENNA__12844__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_180_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_180_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09451_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08402_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ net778 _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08371__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08264_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08226__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12256__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08195_ _03800_ _03805_ net727 vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__mux2_1
XANTENNA__13021__B1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14752__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout405_A _07664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1147_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12272__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1009 net1010 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09623__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout774_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__B2 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ net1078 net1030 net1026 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout941_A _03555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _05325_ _05326_ _05327_ _05328_ net797 net816 vssd1 vssd1 vccd1 vccd1 _05329_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12835__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _06346_ _06477_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__and2_1
X_09649_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__mux2_1
XANTENNA__10310__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14927__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12660_ _07289_ net2526 net475 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09520__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11611_ net574 _07098_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13260__A0 net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08267__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12063__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ _07560_ net482 net412 net2088 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11351__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14330_ net1088 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03489_ _03488_
+ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__a41o_1
XFILLER_0_93_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11542_ _06940_ _07028_ net562 vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\]
+ _03438_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13012__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ net553 _06921_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ clknet_leaf_51_wb_clk_i _01676_ _00229_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_13212_ net90 team_04_WB.MEM_SIZE_REG_REG\[29\] net983 vssd1 vssd1 vccd1 vccd1 _01691_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__07975__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input70_A wbs_dat_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09767__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _03533_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] vssd1 vssd1
+ vccd1 vccd1 _06003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09756__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14192_ _03377_ _03401_ team_04_WB.instance_to_wrap.final_design.v_out vssd1 vssd1
+ vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_state\[0\] sky130_fd_sc_hd__o21a_1
XANTENNA__11574__A0 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ _07577_ net370 net294 net2000 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a22o_1
X_10355_ _05624_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nand2b_1
X_13074_ net256 net2285 net305 vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output157_A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_163_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16902_ clknet_leaf_19_wb_clk_i _02571_ _01131_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\]
+ sky130_fd_sc_hd__dfrtp_1
X_12025_ net258 net684 vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13079__A0 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16833_ clknet_leaf_133_wb_clk_i _02502_ _01062_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16764_ clknet_leaf_127_wb_clk_i _02433_ _00993_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13976_ _04411_ net599 vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__and2b_1
XANTENNA__12826__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15715_ net1295 vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__inv_2
X_12927_ net217 net2279 net318 vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__mux2_1
X_16695_ clknet_leaf_154_wb_clk_i _02364_ _00924_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\]
+ sky130_fd_sc_hd__dfrtp_1
X_15646_ net1180 vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__inv_2
X_12858_ _07558_ net340 net390 net1995 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09430__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11809_ net758 _05830_ net697 _04057_ net693 vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__a221o_1
XANTENNA__12054__B2 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15577_ net1248 vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__inv_2
X_12789_ _07516_ net347 net399 net2319 vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17316_ net1372 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_127_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11261__A _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528_ net1193 vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12076__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17247_ net1307 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_25_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14459_ net1277 vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__inv_2
XANTENNA__12791__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13003__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17178_ clknet_leaf_88_wb_clk_i _02790_ _01407_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10368__B2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16129_ clknet_leaf_136_wb_clk_i _01798_ _00358_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12092__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12109__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__mux2_1
XANTENNA__13857__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_63_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07902_ team_04_WB.instance_to_wrap.final_design.uart.receiving vssd1 vssd1 vccd1
+ vccd1 _03517_ sky130_fd_sc_hd__inv_2
XANTENNA__11868__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08882_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13194__Y _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09605__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13635__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11436__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09503_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout355_A _07484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A1_N net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1097_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09340__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09365_ net627 _04973_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_A _06197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1264_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08316_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\]
+ net929 vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\]
+ net856 vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_41 net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08247_ _03854_ _03855_ _03856_ _03857_ net831 net747 vssd1 vssd1 vccd1 vccd1 _03858_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout310_X net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12348__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ net721 _03788_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout891_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout989_A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10515__A team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _05750_ _05710_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__nand2b_1
Xoutput170 net170 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput181 net181 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput192 net192 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__buf_2
X_10071_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] _04168_ vssd1
+ vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__and2_1
XANTENNA__10802__X _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ _03211_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__nand2_1
XANTENNA__12808__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] net1043 _03151_
+ net1081 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ _04384_ _06460_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_67_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15500_ net1119 vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__inv_2
XANTENNA__10295__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ net2152 net405 net333 _07381_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__a22o_1
X_16480_ clknet_leaf_135_wb_clk_i _02149_ _00709_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13692_ _03068_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14025__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09250__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15431_ net1139 vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__inv_2
XANTENNA__13233__A0 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _07614_ net482 net408 net1786 vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ net1219 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _07541_ net486 net417 net1791 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11795__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17101_ clknet_leaf_104_wb_clk_i _02736_ _01330_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14313_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[17\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[16\] net1091
+ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15488__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11525_ _06910_ _07013_ net563 vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15293_ net1153 vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ clknet_leaf_114_wb_clk_i _02701_ _01261_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
X_14244_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\]
+ _03426_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\] vssd1 vssd1
+ vccd1 vccd1 _03431_ sky130_fd_sc_hd__a31o_1
Xwire275 _07215_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_1
XANTENNA_input73_X net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ _06943_ _06944_ net587 vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10407_ net618 _05988_ net283 vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__a21oi_1
X_14175_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] vssd1 vssd1
+ vccd1 vccd1 _03391_ sky130_fd_sc_hd__and3_1
X_11387_ _04557_ _04584_ net359 _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13126_ _07560_ net377 net296 net1980 vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__a22o_1
X_10338_ _05588_ _05589_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_119_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13057_ _07246_ net2556 net303 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__mux2_1
X_10269_ net621 _05867_ net278 vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09425__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ net2375 net515 _07457_ net440 vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a22o_1
XANTENNA__12511__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11527__Y _07016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_147_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_108_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16816_ clknet_leaf_191_wb_clk_i _02485_ _01045_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[789\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13959_ _03918_ net262 net598 _03313_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a31o_1
X_16747_ clknet_leaf_15_wb_clk_i _02416_ _00976_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13472__B1 team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12275__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16678_ clknet_leaf_22_wb_clk_i _02347_ _00907_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09160__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13224__A0 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13190__B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15629_ net1144 vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17234__1299 vssd1 vssd1 vccd1 vccd1 _17234__1299/HI net1299 sky130_fd_sc_hd__conb_1
XANTENNA__08326__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ net779 _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__nor2_1
XANTENNA__12578__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08101_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08877__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[940\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _03640_ net703 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
XANTENNA__13189__Y _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput61 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_1
XFILLER_0_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11538__B1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput72 wbs_dat_i[12] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_4
Xhold801 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\] vssd1 vssd1
+ vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold812 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\] vssd1 vssd1
+ vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 wbs_dat_i[22] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_1
XFILLER_0_114_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold823 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\] vssd1 vssd1
+ vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_1
XANTENNA__11002__A2 _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold834 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\] vssd1 vssd1
+ vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\] vssd1 vssd1
+ vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\] vssd1 vssd1
+ vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_186_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold867 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\] vssd1 vssd1
+ vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold878 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\] vssd1 vssd1
+ vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 team_04_WB.instance_to_wrap.final_design.uart.working_data\[6\] vssd1 vssd1
+ vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ net629 _04893_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__and2b_1
XANTENNA__10054__B _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1012_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__S net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ net637 _04473_ _04439_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout472_A net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08796_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_154_Right_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout737_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10816__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09070__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13215__A0 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ _05022_ _05027_ net724 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__mux2_1
XANTENNA__12018__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout525_X net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12569__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09348_ net726 _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_134_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ _04886_ _04887_ _04888_ _04889_ net786 net806 vssd1 vssd1 vccd1 vccd1 _04890_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15101__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ net574 _06798_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_151_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12290_ _07443_ _07444_ net675 vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_151_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12444__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11241_ team_04_WB.MEM_SIZE_REG_REG\[19\] _06510_ vssd1 vssd1 vccd1 vccd1 _06730_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_73_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12741__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08945__B2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _03891_ net642 net544 vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _05732_ _05733_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15980_ clknet_leaf_51_wb_clk_i _01656_ _00209_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10054_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _03836_ vssd1
+ vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or2_1
X_14931_ net1231 vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__inv_2
XANTENNA_input33_A DAT_I[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__X _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14862_ net1200 vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__inv_2
X_13813_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] net1043 _03203_
+ net1081 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16601_ clknet_leaf_152_wb_clk_i _02270_ _00830_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_106_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_82_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14793_ net1136 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__inv_2
XANTENNA__12257__B2 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16532_ clknet_leaf_2_wb_clk_i _02201_ _00761_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ net1093 _03134_ net1045 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\]
+ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o2bb2a_1
X_10956_ _06379_ _06427_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__nand3_2
XFILLER_0_35_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16463_ clknet_leaf_187_wb_clk_i _02132_ _00692_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13675_ net1001 _03064_ _03065_ _03063_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10887_ _04723_ _06375_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__and2_1
XFILLER_0_156_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15414_ net1223 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__inv_2
X_12626_ _07597_ net483 net409 net1889 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16394_ clknet_leaf_163_wb_clk_i _02063_ _00623_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15345_ net1271 vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__inv_2
XANTENNA__08633__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12557_ _07524_ net487 net418 net1880 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_171_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13230__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_26 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11508_ _06383_ _06427_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_91_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15276_ net1122 vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12488_ _07485_ net483 net424 net1798 vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a22o_1
XANTENNA__10991__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\] vssd1 vssd1
+ vccd1 vccd1 net1545 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09808__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17015_ clknet_leaf_173_wb_clk_i _02684_ _01244_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\]
+ sky130_fd_sc_hd__dfrtp_1
X_14227_ _07715_ net818 _03420_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__and3_1
Xhold119 _02761_ vssd1 vssd1 vccd1 vccd1 net1556 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ net573 _06831_ _06926_ _06271_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__o211a_1
XANTENNA__14850__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__X _07675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09944__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12732__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ _03373_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13109_ _07541_ net371 net298 net1982 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ net1494 _06124_ net1035 vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__mux2_1
XANTENNA__12496__A1 _07493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1170 net1172 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_4
Xfanout1181 net1187 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__clkbuf_2
X_08650_ net779 _04260_ net761 vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21ai_1
Xfanout1192 net1193 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08994__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__C net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ net716 _04191_ _04180_ _04174_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_87_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10259__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07911__B net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_159_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09202_ net633 net590 vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__nand2_1
XANTENNA__13748__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11208__C1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__mux2_1
XANTENNA__12420__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout220_A _07271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout318_A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__mux2_1
XANTENNA__08234__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08015_ _03625_ _03598_ _03616_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__and3b_1
XANTENNA__10982__B2 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold620 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\] vssd1 vssd1
+ vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\] vssd1 vssd1
+ vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold642 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\] vssd1 vssd1
+ vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold653 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\] vssd1 vssd1
+ vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12723__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__A1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\] vssd1 vssd1
+ vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold675 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1005\] vssd1 vssd1
+ vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\] vssd1 vssd1
+ vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout687_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold697 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\] vssd1 vssd1
+ vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _05575_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ net661 _04526_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__o21ai_4
X_09897_ _03865_ _05507_ net643 _03862_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_A net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08786__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1009\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__mux2_1
X_08779_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ _06291_ _06298_ net658 vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_0_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ net686 _07273_ _07274_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14000__A _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ net636 net550 _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11343__B _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269__1329 vssd1 vssd1 vccd1 vccd1 _17269__1329/HI net1329 sky130_fd_sc_hd__conb_1
XFILLER_0_165_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__X _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13460_ net1002 _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__nand2_1
XANTENNA__10670__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ net1520 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1
+ vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_153_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ net2381 net432 _07633_ net519 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13391_ net1086 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 _07817_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12411__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15130_ net1137 vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__inv_2
X_12342_ net2100 net502 _07615_ net458 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ net1211 vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__inv_2
X_12273_ net2489 net503 _07579_ net441 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14012_ _05307_ _03336_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__nor2_1
X_11224_ _06461_ _06711_ _06459_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12714__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10725__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ net582 _06643_ net288 vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10106_ _04948_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] vssd1
+ vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__and2b_1
XANTENNA_input36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15963_ clknet_leaf_69_wb_clk_i _01639_ _00192_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11086_ _05057_ net551 _06574_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__o21ai_1
X_10037_ _05560_ _05646_ _05562_ _05559_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a211o_1
X_14914_ net1240 vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__inv_2
X_15894_ clknet_leaf_35_wb_clk_i _01571_ _00121_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09703__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14845_ net1149 vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14776_ net1208 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08319__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ net655 _07443_ _07444_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__and3_1
XANTENNA__11989__B1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12349__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ team_04_WB.ADDR_START_VAL_REG\[10\] _03117_ vssd1 vssd1 vccd1 vccd1 _03118_
+ sky130_fd_sc_hd__and2_1
X_16515_ clknet_leaf_122_wb_clk_i _02184_ _00744_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _04920_ _06287_ net657 vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_173_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10661__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ net1000 _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__nor2_1
XANTENNA__09939__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16446_ clknet_leaf_158_wb_clk_i _02115_ _00675_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12609_ _07578_ net482 net412 net2615 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16377_ clknet_leaf_177_wb_clk_i _02046_ _00606_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12402__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10413__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15328_ net1152 vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08082__B2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12084__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15259_ net1114 vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__inv_2
XANTENNA__08989__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12705__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A0 _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13902__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13196__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _05425_ _05430_ net730 vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__mux2_1
Xfanout407 _07664_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout429 _07641_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_129_Left_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09751_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__mux2_1
XANTENNA__12469__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _04309_ _04310_ _04311_ _04312_ net789 net801 vssd1 vssd1 vccd1 vccd1 _04313_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13130__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ _05289_ _05290_ _05291_ _05292_ net835 net746 vssd1 vssd1 vccd1 vccd1 _05293_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07922__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ net751 _03656_ _03726_ net662 vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_146_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15912__Q net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08564_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__mux2_1
XANTENNA__08229__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09193__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[599\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout435_A _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Left_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10652__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13197__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout602_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09116_ net703 _04725_ _04330_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_696 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09047_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__mux2_1
XANTENNA__12157__A0 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08899__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold450 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\] vssd1 vssd1
+ vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10168__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\] vssd1 vssd1
+ vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold472 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\] vssd1 vssd1
+ vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold483 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\] vssd1 vssd1
+ vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold494 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\] vssd1 vssd1
+ vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11380__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__clkbuf_4
Xfanout941 _03555_ vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
X_09949_ net593 _04114_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__or2_1
Xfanout952 net956 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_4
XANTENNA__13657__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout963 net964 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout974 _03548_ vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_2
Xfanout985 _07705_ vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__buf_4
XANTENNA__08759__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13121__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout996 net997 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _07628_ net473 net316 net1609 vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\] vssd1 vssd1
+ vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09523__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11911_ net691 _06915_ _07379_ net614 vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__o211a_4
Xhold1161 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\] vssd1 vssd1
+ vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 net118 vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\] vssd1 vssd1
+ vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_142_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _07593_ net340 net386 net1692 vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\] vssd1 vssd1
+ vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14630_ net1106 vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__inv_2
X_11842_ net613 _07318_ _07319_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__and3_4
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_156_Left_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ net1182 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__inv_2
X_11773_ team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07260_ sky130_fd_sc_hd__a21o_1
XANTENNA__11435__A2 _06923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13512_ _07849_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__xnor2_1
X_16300_ clknet_leaf_107_wb_clk_i _01969_ _00529_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\]
+ sky130_fd_sc_hd__dfrtp_1
X_17280_ net1336 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
X_10724_ _06210_ _06212_ net533 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14492_ net1159 vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__inv_2
X_16231_ clknet_leaf_21_wb_clk_i _01900_ _00460_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\]
+ sky130_fd_sc_hd__dfrtp_1
X_13443_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__inv_2
X_10655_ net1558 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1
+ vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08064__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16162_ clknet_leaf_144_wb_clk_i _01831_ _00391_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\]
+ sky130_fd_sc_hd__dfrtp_1
X_13374_ _07786_ _07787_ _07799_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__o21ba_1
Xclkload17 clknet_leaf_191_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__clkinv_4
X_10586_ _06129_ net1613 net1023 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload28 clknet_leaf_172_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__10417__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output187_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15113_ net1132 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__inv_2
Xclkload39 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload39/X sky130_fd_sc_hd__clkbuf_8
X_12325_ net259 net668 vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__and2_2
X_16093_ clknet_leaf_130_wb_clk_i _01762_ _00322_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12148__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_165_Left_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15044_ net1171 vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__inv_2
X_12256_ _07340_ net675 vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__and2_1
XANTENNA__08602__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11207_ net554 _06606_ _06695_ net568 vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__a211o_1
X_12187_ net245 net648 vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_166_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_166_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _06625_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__nor2_1
X_16995_ clknet_leaf_122_wb_clk_i _02664_ _01224_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11963__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15946_ clknet_leaf_57_wb_clk_i _01623_ _00173_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__dfrtp_1
X_11069_ net640 net549 vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__nand2_1
XANTENNA__12320__B1 _07604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09411__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13657__A1_N net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ clknet_leaf_94_wb_clk_i _01554_ _00104_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\]
+ sky130_fd_sc_hd__dfrtp_4
X_14828_ net1128 vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12794__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14759_ net1137 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08280_ _03872_ _03878_ _03889_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_117_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13179__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ clknet_leaf_43_wb_clk_i _02098_ _00658_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12387__A0 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__B2 team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12139__A0 _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13887__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__C _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_1
Xfanout226 _07289_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__buf_2
XANTENNA__11362__A1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_1
X_09803_ net725 _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__or2_1
XANTENNA__11362__B2 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17268__1328 vssd1 vssd1 vccd1 vccd1 _17268__1328/HI net1328 sky130_fd_sc_hd__conb_1
Xfanout248 _07307_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10062__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] net1077 net1030 net1026 vssd1
+ vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or4_1
Xfanout259 _07349_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_2
XANTENNA_fanout385_A _07674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13103__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09307__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _03507_ net1008 net1007 _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__a32o_1
XANTENNA__14102__X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08748__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09343__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ net768 _05275_ _05264_ _05258_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout552_A _05376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08616_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07964__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ net775 _05200_ _05206_ net763 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__o211a_1
XFILLER_0_167_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09166__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08547_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout817_A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10518__A team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12378__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12436__C net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _06017_ _06018_ _06008_ _06013_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12917__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14119__A1 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14119__B2 team_04_WB.ADDR_START_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11050__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10371_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] _05527_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12292__X _07589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__A3 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ net233 net678 vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09518__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ _07522_ net373 net299 net1924 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a22o_1
XANTENNA__08422__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12041_ net261 net682 vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__and2_2
Xhold280 net145 vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold291 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\] vssd1 vssd1
+ vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout760 _03613_ vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__buf_2
Xfanout771 net777 vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__buf_4
Xfanout782 _03563_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_4
X_16780_ clknet_leaf_111_wb_clk_i _02449_ _01009_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13992_ _04811_ net262 _03325_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__and3_1
Xfanout793 net795 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_161_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_161_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ net1292 vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__inv_2
X_12943_ _07374_ net2557 net321 vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15662_ net1173 vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__inv_2
X_12874_ _07574_ net347 net391 net2560 vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a22o_1
XANTENNA__08945__X _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11825_ team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07305_ sky130_fd_sc_hd__a21o_1
X_14613_ net1200 vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__inv_2
X_15593_ net1132 vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14395__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17332_ net1388 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
X_14544_ net1260 vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11756_ net705 _05777_ net690 _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__o211a_1
XANTENNA__11813__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12081__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _05111_ _06191_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nand2_2
X_17263_ net1323 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_165_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14475_ net1159 vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12369__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ net571 _06226_ _06279_ _07016_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13426_ team_04_WB.MEM_SIZE_REG_REG\[24\] _07736_ _07737_ vssd1 vssd1 vccd1 vccd1
+ _07852_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08037__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12908__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16214_ clknet_leaf_10_wb_clk_i _01883_ _00443_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\]
+ sky130_fd_sc_hd__dfrtp_1
X_17194_ clknet_leaf_79_wb_clk_i _02806_ _01423_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10638_ net1487 net2668 _06173_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload106 clknet_leaf_112_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload106/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload117 clknet_leaf_135_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload128 clknet_leaf_118_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16145_ clknet_leaf_175_wb_clk_i _01814_ _00374_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload139 clknet_leaf_107_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload139/Y sky130_fd_sc_hd__bufinv_16
X_13357_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] team_04_WB.MEM_SIZE_REG_REG\[5\]
+ _07778_ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__and4_1
XANTENNA__09936__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06118_ sky130_fd_sc_hd__and3_1
XANTENNA__10715__X _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_168_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09428__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ net2108 net499 _07598_ net436 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16076_ clknet_leaf_107_wb_clk_i _01745_ _00305_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_13288_ team_04_WB.instance_to_wrap.final_design.uart.receiving _06170_ _07717_ vssd1
+ vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15027_ net1227 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__inv_2
XANTENNA__11259__A net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12239_ net2408 net504 _07562_ net445 vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XANTENNA__08745__C1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16978_ clknet_leaf_9_wb_clk_i _02647_ _01207_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput4 DAT_I[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09163__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15929_ clknet_leaf_59_wb_clk_i _01606_ _00156_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08401_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09381_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\]
+ net951 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _03939_ _03940_ _03941_ _03942_ net788 net809 vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08371__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_717 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08263_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\]
+ net930 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_92_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08194_ _03801_ _03802_ _03803_ _03804_ net826 net750 vssd1 vssd1 vccd1 vccd1 _03805_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10057__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12780__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_669 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12272__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09528__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09623__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout767_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13384__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ net765 _03588_ _03577_ _03576_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__09073__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\]
+ net970 vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__mux2_1
XANTENNA__11616__B _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_X net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09139__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ _05184_ _05189_ net724 vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12599__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ net568 _06911_ _06278_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__a21o_1
XANTENNA__15104__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__A1 team_04_WB.ADDR_START_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12590_ _07559_ net487 net414 net2134 vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a22o_1
XANTENNA__12063__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11351__B _06839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ net568 _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\]
+ _03437_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\] vssd1 vssd1
+ vccd1 vccd1 _03441_ sky130_fd_sc_hd__a31o_1
XFILLER_0_163_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13012__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ net539 _06583_ _06585_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__nand3_1
XFILLER_0_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13211_ net92 team_04_WB.MEM_SIZE_REG_REG\[30\] net982 vssd1 vssd1 vccd1 vccd1 _01692_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03528_
+ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_1
X_14191_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\] _03400_
+ _03373_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_115_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11574__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12771__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09248__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13142_ _07576_ net371 net295 net2368 vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a22o_1
XANTENNA_input63_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nor2_1
XANTENNA__08152__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11079__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _07356_ net2403 net304 vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__mux2_1
X_10285_ _05573_ _05574_ _05637_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_163_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16901_ clknet_leaf_170_wb_clk_i _02570_ _01130_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\]
+ sky130_fd_sc_hd__dfrtp_1
X_12024_ net2397 net516 _07465_ net446 vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_163_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_168_Right_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11877__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__S1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_137_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16832_ clknet_leaf_138_wb_clk_i _02501_ _01061_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11807__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16763_ clknet_leaf_100_wb_clk_i _02432_ _00992_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\]
+ sky130_fd_sc_hd__dfrtp_1
X_13975_ _04355_ net263 net598 _03321_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15714_ net1261 vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__inv_2
X_12926_ net220 net2434 net320 vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__mux2_1
X_16694_ clknet_leaf_12_wb_clk_i _02363_ _00923_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11813__Y _07295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15645_ net1180 vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__inv_2
X_12857_ _07557_ net334 net389 net2118 vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13233__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11808_ net2436 net526 net438 _07290_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15576_ net1221 vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__inv_2
X_12788_ _07515_ net344 net398 net1817 vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XANTENNA__12054__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12357__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17315_ net1371 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
X_14527_ net1193 vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__inv_2
X_11739_ _06918_ _06957_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17267__1327 vssd1 vssd1 vccd1 vccd1 _17267__1327/HI net1327 sky130_fd_sc_hd__conb_1
XFILLER_0_3_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11801__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17246_ net1306 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XANTENNA__09947__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13003__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14458_ net1278 vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ _07827_ _07834_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__nor2_1
XANTENNA__10592__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17177_ clknet_leaf_88_wb_clk_i _02789_ _01406_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_14389_ net1466 vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09158__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12762__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16128_ clknet_leaf_140_wb_clk_i _01797_ _00357_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_176_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12092__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux2_1
X_16059_ clknet_leaf_104_wb_clk_i _01728_ _00288_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12514__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ net1 vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__inv_2
X_08881_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1008\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_102_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13635__C net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09502_ _03643_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or2_2
XFILLER_0_154_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09621__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09433_ net774 _05037_ net763 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout348_A net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ net627 _04973_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_164_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08249__B2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_111_Left_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08315_ net773 _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09295_ net728 _04905_ net712 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__o21a_1
XANTENNA_31 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout515_A _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1257_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\]
+ net883 vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13488__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _03784_ _03785_ _03786_ _03787_ net826 net742 vssd1 vssd1 vccd1 vccd1 _03788_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A1 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12753__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09068__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10515__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_A net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput160 net160 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput171 net171 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_120_Left_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12505__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput182 net182 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput193 net193 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
X_10070_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _04113_ vssd1
+ vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nand2_1
XANTENNA__11859__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08700__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11627__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ _07834_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ _04385_ _06460_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12711_ net2280 net405 net338 _07375_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13691_ _03079_ _03080_ _03074_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09780__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__A net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15430_ net1103 vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__inv_2
X_12642_ _07613_ net479 net408 net1851 vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12036__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12177__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ net1167 vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_156_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _07540_ net488 net418 net1780 vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_363 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11795__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17100_ clknet_leaf_105_wb_clk_i _02735_ _01329_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14312_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[29\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[28\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[25\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[24\] net1090
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\] vssd1 vssd1
+ vccd1 vccd1 _03472_ sky130_fd_sc_hd__mux4_1
XANTENNA__11795__B2 net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ net630 net628 net627 net589 net546 net540 vssd1 vssd1 vccd1 vccd1 _07013_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15292_ net1148 vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14243_ net2657 _03428_ _03430_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17031_ clknet_leaf_165_wb_clk_i _02700_ _01260_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
X_11455_ net562 _06240_ _06571_ _06937_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__a31o_1
Xwire276 _07210_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12193__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12744__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1059 vssd1
+ vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__xnor2_1
X_14174_ _03389_ _03390_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ _04557_ _04584_ net360 vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ _07559_ net376 net296 net1925 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a22o_1
X_10337_ _05750_ _05927_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13056_ _07657_ _07666_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__or2_4
X_10268_ _05760_ _05761_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08610__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13228__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ net241 net680 vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__and2_1
XANTENNA__15009__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _05651_ _05804_ _05805_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_159_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_159_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16815_ clknet_leaf_189_wb_clk_i _02484_ _01044_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14848__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16746_ clknet_leaf_166_wb_clk_i _02415_ _00975_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12275__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ net155 net1064 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__and2_1
XANTENNA__09441__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _07611_ net339 net385 net1927 vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16677_ clknet_leaf_4_wb_clk_i _02346_ _00906_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\]
+ sky130_fd_sc_hd__dfrtp_1
X_13889_ _03258_ _03268_ net2623 net1066 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_159_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15628_ net1119 vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__inv_2
XANTENNA__13224__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__A1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08326__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ net1141 vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15791__10 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__inv_2
X_08100_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12983__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09080_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1004\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08031_ _03591_ net759 net752 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput40 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13199__A _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17229_ net1435 _02839_ _01485_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput51 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold802 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\] vssd1 vssd1
+ vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
Xinput62 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_102_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput73 wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_1
XANTENNA__12735__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput84 wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_1
Xhold813 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\] vssd1 vssd1
+ vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 wbs_dat_i[4] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__buf_1
XFILLER_0_141_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold824 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\] vssd1 vssd1
+ vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\] vssd1 vssd1
+ vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\] vssd1 vssd1
+ vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10210__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold857 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\] vssd1 vssd1
+ vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09982_ _04893_ net628 vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__and2b_1
Xhold868 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\] vssd1 vssd1
+ vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold879 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\] vssd1 vssd1
+ vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_61 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09616__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08933_ net781 _04543_ net764 vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15915__Q net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13160__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _04439_ net637 _04473_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__or3_1
XFILLER_0_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10070__B _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout465_A _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14110__X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout253_X net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout632_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09416_ _05023_ _05024_ _05025_ _05026_ net831 net747 vssd1 vssd1 vccd1 vccd1 _05027_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_95_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12018__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10029__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11226__A0 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09347_ _04954_ _04955_ _04956_ _04957_ net836 net748 vssd1 vssd1 vccd1 vccd1 _04958_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_165_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11777__A1 _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12974__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11529__A1 _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12444__C net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12726__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ net463 _06712_ _06713_ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o31a_1
XFILLER_0_160_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _06658_ _06659_ net463 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10122_ net1059 _05283_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__or2_1
XANTENNA__08430__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__and2b_1
X_14930_ net1238 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266__1326 vssd1 vssd1 vccd1 vccd1 _17266__1326/HI net1326 sky130_fd_sc_hd__conb_1
XANTENNA__14326__S0 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A DAT_I[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ net1210 vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14100__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ clknet_leaf_149_wb_clk_i _02269_ _00829_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\]
+ sky130_fd_sc_hd__dfrtp_1
X_13812_ _07854_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_106_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14792_ net1124 vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__inv_2
XANTENNA__12257__A2 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16531_ clknet_leaf_182_wb_clk_i _02200_ _00760_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[504\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13743_ _07777_ _07803_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_158_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10955_ _06383_ _06437_ _06443_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_27_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16462_ clknet_leaf_27_wb_clk_i _02131_ _00691_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[435\]
+ sky130_fd_sc_hd__dfrtp_1
X_13674_ net1098 _03061_ net1046 net1059 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13206__B2 team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10886_ _04753_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15413_ net1214 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _07596_ net485 net409 net1728 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a22o_1
X_16393_ clknet_leaf_101_wb_clk_i _02062_ _00622_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11768__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12965__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12556_ _07523_ net481 net416 net1835 vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a22o_1
X_15344_ net1162 vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _06503_ _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12127__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12980__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ net1122 vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__inv_2
X_12487_ net699 _06198_ _07483_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__or3_4
XFILLER_0_110_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12717__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold109 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[14\] vssd1
+ vssd1 vccd1 vccd1 net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17014_ clknet_leaf_14_wb_clk_i _02683_ _01243_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\]
+ sky130_fd_sc_hd__dfrtp_1
X_14226_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11438_ _04530_ net363 net362 _04529_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14157_ _03527_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__and2_1
XANTENNA__13747__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11369_ net706 _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__nor2_1
XANTENNA__09944__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13108_ _07540_ net380 net301 net1677 vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a22o_1
X_14088_ net1500 _06122_ net1033 vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__mux2_1
XANTENNA__08340__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13142__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13039_ _07500_ net375 net307 net1714 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a22o_1
XANTENNA__12496__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09897__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1166 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09960__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_4
XANTENNA__14317__S0 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1182 net1183 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
XANTENNA__12797__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14578__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13482__A team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08580_ _04185_ _04190_ net721 vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1003 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10259__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16729_ clknet_leaf_152_wb_clk_i _02398_ _00958_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11456__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12098__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08321__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09201_ _03628_ _03644_ _04811_ net666 _04780_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__a221oi_4
Xclkbuf_leaf_56_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09132_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12420__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[492\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[460\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout213_A _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ _03600_ _03602_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__or4_1
XANTENNA__12708__B1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold610 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\] vssd1 vssd1
+ vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold621 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\] vssd1 vssd1
+ vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10065__B _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\] vssd1 vssd1
+ vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\] vssd1 vssd1
+ vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12184__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10853__A_N _04166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\] vssd1 vssd1
+ vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09854__B net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14105__X net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold665 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\] vssd1 vssd1
+ vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\] vssd1 vssd1
+ vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1122_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold687 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\] vssd1 vssd1
+ vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08250__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\] vssd1 vssd1
+ vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand2_1
XANTENNA__12280__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _03558_ net702 _04386_ net662 vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__a211o_1
X_09896_ _03781_ _03808_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__nor2_1
XANTENNA__10512__C net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08786__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _04451_ _04452_ _04457_ net731 net715 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__mux2_1
XANTENNA__12239__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13987__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout635_X net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14000__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ net665 _05375_ _05340_ _04440_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_101_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10670__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_10671_ net2648 net1018 net1014 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1
+ vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12947__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ net651 net600 net237 vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_11_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13390_ _07768_ _07815_ _07764_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12411__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ net249 net671 vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12962__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15060_ net1235 vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__inv_2
X_12272_ net251 net672 vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14011_ net1642 net1069 _03341_ net264 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a22o_1
XANTENNA__13567__A team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _06459_ _06461_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11922__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ net571 _06642_ _06532_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__a21o_1
XANTENNA__13124__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _04893_ vssd1
+ vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nand2_1
X_15962_ clknet_leaf_71_wb_clk_i _01638_ _00191_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11085_ net580 net551 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__nand2_1
XANTENNA__13675__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ _05560_ _05646_ _05562_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__a21o_1
X_14913_ net1150 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output132_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ clknet_leaf_30_wb_clk_i _01570_ _00120_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11150__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ net1126 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11438__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14775_ net1226 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ _07443_ _07444_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__and2_2
XFILLER_0_169_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16514_ clknet_leaf_146_wb_clk_i _02183_ _00743_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\]
+ sky130_fd_sc_hd__dfrtp_1
X_13726_ _07696_ _03111_ _03113_ net999 _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10938_ _06392_ _06396_ _06422_ _06426_ _06425_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__a41o_2
XANTENNA__12650__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16445_ clknet_leaf_129_wb_clk_i _02114_ _00674_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\]
+ sky130_fd_sc_hd__dfrtp_1
X_13657_ net1098 _03047_ net1046 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09939__B _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ _06286_ _06289_ _06293_ _05463_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__a31o_1
XANTENNA__10661__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10718__X _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12938__A0 _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13241__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11550__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _07577_ net485 net413 net2107 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16376_ clknet_leaf_149_wb_clk_i _02045_ _00605_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12402__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ team_04_WB.ADDR_START_VAL_REG\[13\] _02971_ _02975_ _02978_ vssd1 vssd1 vccd1
+ vccd1 _02979_ sky130_fd_sc_hd__and4_1
XFILLER_0_155_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10413__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15327_ net1249 vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12539_ net2130 net256 net423 vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_87 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15258_ net1138 vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14209_ net1087 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ _03409_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14072__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A1 _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15189_ net1207 vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_174_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_174_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13196__B net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _07661_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout419 _07659_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_103_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13115__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _05349_ _05355_ _05360_ net732 net715 vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__o221a_1
XANTENNA__12469__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\]
+ net937 vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08632_ _04225_ _04231_ _04242_ net716 vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a22o_4
XANTENNA__07922__B net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13825__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ net721 _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11524__S0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08494_ _04101_ _04102_ _04103_ _04104_ net784 net805 vssd1 vssd1 vccd1 vccd1 _04105_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09193__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12641__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10652__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1072_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A _07641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08245__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17265__1325 vssd1 vssd1 vccd1 vccd1 _17265__1325/HI net1325 sky130_fd_sc_hd__conb_1
XFILLER_0_134_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09115_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout797_A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold440 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\] vssd1 vssd1
+ vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold451 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\] vssd1
+ vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__A1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\] vssd1 vssd1
+ vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09076__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold473 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\] vssd1 vssd1
+ vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold484 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\] vssd1 vssd1
+ vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold495 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\] vssd1 vssd1
+ vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout920 net926 vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__buf_2
XANTENNA__13106__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 net941 vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09948_ net596 _04056_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__xnor2_1
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout953 net956 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout964 net972 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_4
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09804__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout986 net988 vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08759__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout997 net998 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _04923_ _04947_ _04974_ _04920_ net629 vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\] vssd1 vssd1
+ vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\] vssd1 vssd1
+ vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net688 _07376_ _07378_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__a21o_1
XANTENNA__15107__A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1162 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\] vssd1 vssd1
+ vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\] vssd1 vssd1
+ vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12890_ _07592_ net335 net385 net2376 vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\] vssd1 vssd1
+ vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12880__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1195 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\] vssd1 vssd1
+ vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_246 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11841_ _06786_ _06815_ net689 vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_16_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14946__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14560_ net1184 vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ net1907 net528 net440 _07259_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XANTENNA__11073__C _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12632__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13511_ _07742_ _07846_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__nor2_1
X_10723_ _05336_ net552 _06211_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__a21o_1
XFILLER_0_126_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14491_ net1120 vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13061__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16230_ clknet_leaf_19_wb_clk_i _01899_ _00459_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input93_A wbs_dat_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13442_ team_04_WB.MEM_SIZE_REG_REG\[28\] _07860_ _07867_ vssd1 vssd1 vccd1 vccd1
+ _07868_ sky130_fd_sc_hd__a21o_1
X_10654_ net1623 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1
+ vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__a22o_1
XANTENNA__12185__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13373_ _07792_ _07798_ _07788_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__o21a_1
X_16161_ clknet_leaf_141_wb_clk_i _01830_ _00390_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[5\]
+ _06128_ net1050 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__mux2_1
Xclkload18 clknet_leaf_192_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__14681__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload29 clknet_leaf_174_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
X_15112_ net1118 vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09775__A net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ net2345 net502 _07606_ net459 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_1_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16092_ clknet_leaf_128_wb_clk_i _01761_ _00321_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_15043_ net1165 vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__inv_2
X_12255_ net2483 net504 _07570_ net447 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12699__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11206_ net554 _06594_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__nor2_1
X_12186_ net2009 net508 _07534_ net447 vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_166_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ team_04_WB.MEM_SIZE_REG_REG\[29\] _06517_ vssd1 vssd1 vccd1 vccd1 _06626_
+ sky130_fd_sc_hd__xor2_2
X_16994_ clknet_leaf_139_wb_clk_i _02663_ _01223_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09714__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15945_ clknet_leaf_57_wb_clk_i _01622_ _00172_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__dfrtp_1
X_11068_ net595 net543 _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13236__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _05587_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__nor2_1
XANTENNA__12140__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ clknet_leaf_94_wb_clk_i _01553_ _00103_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12871__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14827_ net1168 vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14758_ net1111 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__inv_2
XANTENNA__12623__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13709_ _07769_ _07813_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__xor2_1
XANTENNA__10595__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14067__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14689_ net1148 vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__inv_2
XFILLER_0_172_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ clknet_leaf_107_wb_clk_i _02097_ _00657_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_82_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10608__B _06145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15687__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16359_ clknet_leaf_165_wb_clk_i _02028_ _00588_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08686__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14128__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09802_ _05409_ _05410_ _05411_ _05412_ net834 net738 vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__mux4_1
Xfanout227 _07283_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
X_07994_ net1080 net1029 net1025 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a31o_1
Xfanout249 net250 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
XFILLER_0_158_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ net1008 net1007 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\]
+ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09851__C _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08515__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09664_ _05269_ _05274_ net775 vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__mux2_1
XANTENNA__12862__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08615_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[244\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
X_09595_ net780 _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_71_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_173_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1287_A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08546_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__mux2_1
XANTENNA__09166__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11822__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08913__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ _03920_ _03977_ _04031_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__and4_1
XANTENNA__12286__A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout712_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10518__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_196 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11050__A1 _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14119__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_149_Right_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ net1057 _05953_ _05956_ _05957_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_60_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ _04634_ _04639_ net726 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__mux2_1
XANTENNA__14006__A _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_148_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12452__C net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ net2503 net518 _07473_ net458 vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
Xhold270 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\] vssd1 vssd1
+ vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\] vssd1 vssd1
+ vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\] vssd1 vssd1
+ vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11917__X _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__A1 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_144_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_127_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout750 _03648_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09534__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout761 _03570_ vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_8
Xfanout772 net773 vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
Xfanout783 net790 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__clkbuf_8
X_13991_ net1442 net1064 _03330_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a21o_1
Xfanout794 net795 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__buf_4
X_15730_ net1292 vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_161_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _07368_ net2498 net320 vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_161_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08010__Y _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15661_ net1173 vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_2
X_12873_ _07573_ net350 net390 net2095 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a22o_1
XANTENNA__14055__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14612_ net1208 vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__inv_2
X_11824_ net758 _05845_ net697 _04168_ net693 vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__a221o_1
X_15592_ net1116 vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__inv_2
XANTENNA__12605__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17331_ net1387 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_139_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14543_ net1260 vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__inv_2
X_11755_ net686 _07242_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17262_ net1322 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XFILLER_0_154_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ net701 _06183_ _06194_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__or3_4
XANTENNA_input96_X net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ net1273 vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__inv_2
X_11686_ net289 _07171_ _07173_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16213_ clknet_leaf_33_wb_clk_i _01882_ _00442_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\]
+ sky130_fd_sc_hd__dfrtp_1
X_13425_ _07739_ _07846_ _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a21oi_1
X_17193_ clknet_leaf_80_wb_clk_i _02805_ _01422_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net1541 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\] _06173_
+ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13030__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload107 clknet_leaf_113_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload107/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload118 clknet_leaf_136_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15300__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16144_ clknet_leaf_0_wb_clk_i _01813_ _00373_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload129 clknet_leaf_124_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__09709__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13356_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] team_04_WB.MEM_SIZE_REG_REG\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10568_ _06117_ net1553 net1021 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_166_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_168_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11592__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ _07289_ net668 vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__and2_1
XANTENNA__12135__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16075_ clknet_leaf_22_wb_clk_i _01744_ _00304_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_10499_ _06044_ _06052_ _06054_ _06071_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__a31o_1
X_13287_ _06169_ _07713_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_15_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ net1238 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__inv_2
X_12238_ net227 net673 vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__and2_1
XANTENNA__09093__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__A1 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__X _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ net217 net648 vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__and2_1
XANTENNA__09444__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16977_ clknet_leaf_180_wb_clk_i _02646_ _01206_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13097__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput5 DAT_I[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_17264__1324 vssd1 vssd1 vccd1 vccd1 _17264__1324/HI net1324 sky130_fd_sc_hd__conb_1
X_15928_ clknet_leaf_70_wb_clk_i _01605_ _00155_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12844__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15859_ clknet_leaf_98_wb_clk_i _01536_ _00086_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_149_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14046__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08400_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09380_ net774 _04984_ _04990_ net763 vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08331_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__A1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08262_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\]
+ net930 vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__mux2_1
XANTENNA__07909__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08193_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[956\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__mux2_1
XANTENNA__13021__A2 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09619__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07928__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09528__A2 _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10073__B _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12532__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _03582_ _03587_ net772 vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13952__X _03310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[992\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__mux2_1
XANTENNA__12835__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ net775 _05257_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nor2_1
XFILLER_0_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14037__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09139__S1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ _05185_ _05186_ _05187_ _05188_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05189_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08529_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11540_ _06738_ _06939_ net561 vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ net539 _06938_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ net93 team_04_WB.MEM_SIZE_REG_REG\[31\] net982 vssd1 vssd1 vccd1 vccd1 _01693_
+ sky130_fd_sc_hd__mux2_1
X_10422_ _03513_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__or2_1
XANTENNA__09767__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] _03371_
+ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08433__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11574__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\] net1057 _05939_
+ _05942_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a22o_1
X_13141_ _07575_ net380 net296 net2412 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13072_ net259 net2420 net303 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
XANTENNA_input56_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _05573_ _05574_ _05637_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__or3_1
XANTENNA__12523__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16900_ clknet_leaf_173_wb_clk_i _02569_ _01129_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\]
+ sky130_fd_sc_hd__dfrtp_1
X_12023_ net259 net685 vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_163_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09264__S net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ clknet_leaf_159_wb_clk_i _02500_ _01060_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11807__B net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__B _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _05166_ vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_2
XANTENNA__09378__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16762_ clknet_leaf_37_wb_clk_i _02431_ _00991_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\]
+ sky130_fd_sc_hd__dfrtp_1
X_13974_ net146 net1065 vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__and2_1
XANTENNA__12826__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15713_ net1264 vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__inv_2
X_12925_ net214 net2418 net320 vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__mux2_1
X_16693_ clknet_leaf_13_wb_clk_i _02362_ _00922_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[666\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11823__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15644_ net1177 vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12856_ net701 _07555_ _07663_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__or3_4
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ net651 net226 vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15575_ net1231 vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__inv_2
X_12787_ _07514_ net344 net398 net1843 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17314_ net1370 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12357__C net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ net1193 vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11738_ _07151_ _07152_ _07226_ _06841_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__o211a_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11969__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17245_ net1305 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
X_14457_ net1292 vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__inv_2
X_11669_ net530 _06559_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ team_04_WB.MEM_SIZE_REG_REG\[19\] _07746_ _07833_ vssd1 vssd1 vccd1 vccd1
+ _07834_ sky130_fd_sc_hd__a21o_1
XANTENNA__09439__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17176_ clknet_leaf_90_wb_clk_i _02788_ _01405_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_14388_ net1470 vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11565__A2 _06923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ clknet_leaf_154_wb_clk_i _01796_ _00356_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_13339_ net1086 team_04_WB.MEM_SIZE_REG_REG\[12\] vssd1 vssd1 vccd1 vccd1 _07765_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10605__C net47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16058_ clknet_leaf_44_wb_clk_i _01727_ _00287_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07900_ net1092 vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__inv_2
X_15009_ net1188 vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__inv_2
XANTENNA__14080__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08880_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\]
+ net930 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__mux2_1
XANTENNA__10902__A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08813__S0 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10289__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ net719 _03722_ _05111_ _03637_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__a22o_1
XANTENNA__14019__A1 _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07930__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ net780 _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09203__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _04973_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout243_A _07374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ _03921_ _03922_ _03923_ _03924_ net787 net810 vssd1 vssd1 vccd1 vccd1 _03925_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_23_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _04901_ _04902_ _04903_ _04904_ net826 net734 vssd1 vssd1 vccd1 vccd1 _04905_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12450__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _07692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08245_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\]
+ net878 vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__mux2_1
XANTENNA_43 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout410_A _07661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14108__X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout508_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08176_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\]
+ net857 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10515__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput150 net150 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput161 net161 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xoutput172 net172 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__A _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput183 net183 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput194 net194 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__buf_2
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11627__B _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_X net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09812__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _04412_ _06455_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12710_ net2104 net407 net346 _07369_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13690_ _03079_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__nand2_1
XANTENNA__08428__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09113__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _07612_ net486 net408 net2013 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15360_ net1212 vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__inv_2
X_12572_ _07539_ net492 net419 net1711 vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XANTENNA__12441__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14311_ net1090 _03519_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__and2_1
X_11523_ _06424_ _06426_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15291_ net1114 vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17030_ clknet_leaf_19_wb_clk_i _02699_ _01259_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14242_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] _03428_ net819
+ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08163__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11454_ net577 _06941_ _06942_ _06251_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__a211oi_1
X_17263__1323 vssd1 vssd1 vccd1 vccd1 _17263__1323/HI net1323 sky130_fd_sc_hd__conb_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12193__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _05731_ _05740_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__xor2_1
X_14173_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _03387_
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11385_ _06228_ _06669_ _06873_ net585 vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13124_ _07558_ net376 net296 net2078 vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10336_ _05709_ _05710_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10267_ _05569_ _05570_ _05640_ net620 vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o31a_1
X_13055_ _07516_ net383 net309 net1616 vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__a22o_1
XANTENNA__08399__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ net2249 net515 _07456_ net438 vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__a22o_1
X_10198_ _05651_ _05804_ net621 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__o21ai_1
X_16814_ clknet_leaf_42_wb_clk_i _02483_ _01043_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09722__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16745_ clknet_leaf_122_wb_clk_i _02414_ _00974_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\]
+ sky130_fd_sc_hd__dfrtp_1
X_13957_ net1543 net1069 _03312_ net264 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09220__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11483__A1 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12680__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _07610_ net346 net386 net1902 vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__a22o_1
XANTENNA__11483__B2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16676_ clknet_leaf_170_wb_clk_i _02345_ _00905_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\]
+ sky130_fd_sc_hd__dfrtp_1
X_13888_ _02943_ _03194_ _03198_ _03243_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_128_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15627_ net1159 vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12839_ _07537_ net338 net392 net2050 vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a22o_1
XANTENNA__14864__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15558_ net1103 vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08862__A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14509_ net1259 vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14075__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ net1131 vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08030_ _03591_ net759 net752 vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17228_ net1434 _02838_ _01483_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput30 DAT_I[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08073__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput41 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput52 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput63 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold803 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\] vssd1 vssd1
+ vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 wbs_dat_i[14] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_1
X_17159_ clknet_leaf_77_wb_clk_i _02771_ _01388_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold814 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\] vssd1 vssd1
+ vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 wbs_dat_i[24] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_1
Xhold825 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\] vssd1 vssd1
+ vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xinput96 wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_123_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold836 team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\] vssd1 vssd1
+ vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold847 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\] vssd1 vssd1
+ vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold858 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[875\] vssd1 vssd1
+ vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09981_ _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__nand2_1
Xhold869 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[403\] vssd1 vssd1
+ vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08801__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11287__X _06776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _04539_ _04540_ _04541_ _04542_ net798 net803 vssd1 vssd1 vccd1 vccd1 _04543_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12499__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08863_ net637 _04473_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__or2_1
XANTENNA__11171__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08794_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__mux2_1
XANTENNA__09632__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09869__A1_N net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout458_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12671__A0 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08248__S net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12278__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09419__A1 _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10029__A2 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09346_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[424\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\]
+ net899 vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
XANTENNA__09868__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11777__A2 _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__A1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10807__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08228_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__mux2_1
X_11170_ _06352_ _06657_ _06478_ _06345_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__o211ai_1
XANTENNA__09807__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net1059 _05283_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10542__A team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14014__A _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _03493_ _03728_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__nand2_1
XANTENNA__11162__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13853__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16002__Q team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ net1128 vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__inv_2
XANTENNA__14326__S1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14100__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13811_ _07734_ _07737_ _07853_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__and3_1
XANTENNA_input19_A DAT_I[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ net1137 vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13064__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16530_ clknet_leaf_9_wb_clk_i _02199_ _00759_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13742_ _07009_ net271 net710 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10954_ _06442_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__inv_2
XANTENNA__11465__B2 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16461_ clknet_leaf_40_wb_clk_i _02130_ _00690_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ _07090_ net271 _06174_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10885_ _04697_ _06286_ _06294_ net659 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ net1237 vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12624_ _07595_ net482 net408 net1584 vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16392_ clknet_leaf_118_wb_clk_i _02061_ _00621_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12414__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15343_ net1199 vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12555_ _07522_ net483 net417 net2028 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08633__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10717__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ team_04_WB.MEM_SIZE_REG_REG\[8\] _06502_ vssd1 vssd1 vccd1 vccd1 _06995_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15274_ net1106 vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12486_ net2453 net431 net492 _07481_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17013_ clknet_leaf_35_wb_clk_i _02682_ _01242_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\]
+ sky130_fd_sc_hd__dfrtp_1
X_14225_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\] net818 vssd1
+ vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11437_ net573 _06826_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09717__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ _03374_ _03375_ _03530_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11368_ _06842_ _06843_ _06856_ net287 vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__08621__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13239__S net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ _07539_ net382 net301 net1683 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a22o_1
XANTENNA__11548__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10319_ _05908_ _05912_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\]
+ net1056 vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ net1482 _06120_ net1033 vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__mux2_1
X_11299_ net541 _06570_ _06787_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__o21ai_1
X_13038_ _07499_ net382 net309 net1879 vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1150 net1156 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__buf_2
XANTENNA__09960__B _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1161 net1166 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_4
XANTENNA__14317__S1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1172 net1187 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__clkbuf_4
Xfanout1183 net1187 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__buf_4
Xfanout1194 net35 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09452__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14989_ net1152 vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16728_ clknet_leaf_149_wb_clk_i _02397_ _00957_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12098__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08321__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ clknet_leaf_183_wb_clk_i _02328_ _00888_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09200_ _04793_ _04799_ _04810_ net716 vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a22o_4
XFILLER_0_119_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09131_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10967__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09821__B2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09062_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[300\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_96_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_7_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08013_ _03604_ _03618_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold600 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\] vssd1 vssd1
+ vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold611 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\] vssd1 vssd1
+ vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold622 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\] vssd1 vssd1
+ vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12184__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold633 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\] vssd1 vssd1
+ vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09627__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07936__A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold644 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\] vssd1 vssd1
+ vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold655 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\] vssd1 vssd1
+ vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\] vssd1 vssd1
+ vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\] vssd1 vssd1
+ vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold688 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\] vssd1 vssd1
+ vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09964_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__or2_1
Xhold699 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\] vssd1 vssd1
+ vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1115_A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08915_ _04508_ _04514_ _04525_ net716 vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a22o_4
XANTENNA__10081__B _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _04142_ _04194_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__and3b_1
XANTENNA__14769__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__X _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10498__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _04453_ _04454_ _04455_ _04456_ net837 net740 vssd1 vssd1 vccd1 vccd1 _04457_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14121__X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12892__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__S net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__B net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout742_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262__1322 vssd1 vssd1 vccd1 vccd1 _17262__1322/HI net1322 sky130_fd_sc_hd__conb_1
XFILLER_0_67_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12644__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11998__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10670_ net1640 net1018 net1014 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1
+ vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a22o_1
XANTENNA__10670__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09329_ _04936_ _04937_ _04938_ _04939_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04940_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_166 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12340_ net2139 net499 _07614_ net441 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ net2570 net503 _07578_ net442 vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14010_ _05248_ _03336_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__nor2_1
X_11222_ _06454_ _06471_ _06466_ _06462_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_120_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09537__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08441__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13059__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ net554 _06641_ _06534_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_102_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10104_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__inv_2
X_15961_ clknet_leaf_71_wb_clk_i _01637_ _00190_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11084_ net588 net579 net551 vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__mux2_1
XANTENNA__09879__B2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ net592 _04167_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__o21a_1
X_14912_ net1217 vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__inv_2
XANTENNA__10489__A2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12883__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15892_ clknet_leaf_35_wb_clk_i _01569_ _00119_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ net1124 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__inv_2
XANTENNA__12199__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ net1225 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__inv_2
XANTENNA__12635__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ net692 _07057_ net614 vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__o21a_2
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11989__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16513_ clknet_leaf_130_wb_clk_i _02182_ _00742_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ net999 _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _06386_ _06387_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16444_ clknet_leaf_116_wb_clk_i _02113_ _00673_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13656_ _07794_ _07795_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10661__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ net636 _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13060__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ _07576_ net486 net413 net2044 vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16375_ clknet_leaf_167_wb_clk_i _02044_ _00604_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\]
+ sky130_fd_sc_hd__dfrtp_1
X_13587_ net1002 _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12138__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10799_ net590 _04865_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15326_ net1215 vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ net2173 net258 net423 vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11977__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_66 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15257_ net1246 vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12469_ net521 net605 _07470_ net429 net1756 vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a32o_1
X_14208_ net1888 _03409_ _03411_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12166__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net1227 vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__inv_2
XANTENNA__08351__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ net1089 _03361_ net1087 net1088 vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout409 _07661_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09971__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13493__A team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__mux2_1
XANTENNA__12874__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10910__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08631_ _04236_ _04241_ net720 vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ _04169_ _04170_ _04171_ _04172_ net825 net734 vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12626__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08493_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10652__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08526__S net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13051__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout323_A _07671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_A _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09114_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[13\] team_04_WB.instance_to_wrap.CPU_DAT_O\[13\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__mux2_4
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09993__A_N net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09045_ net773 _04649_ net762 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07937__Y _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09357__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11459__Y _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\] vssd1 vssd1
+ vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08114__X _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold441 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\] vssd1 vssd1
+ vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold452 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\] vssd1 vssd1
+ vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 net130 vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11904__A2 _06972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold474 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\] vssd1 vssd1
+ vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold485 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\] vssd1 vssd1
+ vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\] vssd1 vssd1
+ vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_117_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout910 net926 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_2
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09947_ net641 _04003_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2_1
Xfanout932 net934 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__clkbuf_4
Xfanout943 net950 vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
XANTENNA_fanout480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14499__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 net956 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout965 net966 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
Xfanout976 net978 vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_4
X_15807__26 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__inv_2
XANTENNA__10820__A net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _04586_ _04610_ _04643_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a31oi_1
XANTENNA__12865__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout998 _07686_ vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__buf_2
Xhold1130 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\] vssd1 vssd1
+ vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 net171 vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09092__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\] vssd1 vssd1
+ vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ net768 _04432_ _04438_ _04425_ _04426_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__a32o_4
Xhold1163 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\] vssd1 vssd1
+ vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1174 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[385\] vssd1 vssd1
+ vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1185 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\] vssd1 vssd1
+ vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\] vssd1 vssd1
+ vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ net686 _07317_ _07316_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__a21o_1
XANTENNA__12617__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ net653 net212 vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ _07183_ net272 net709 vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10722_ net551 _05404_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nor2_1
XANTENNA__11840__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08436__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490_ net1120 vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_172_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _07726_ _07866_ _07860_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__o21ba_1
X_10653_ net1573 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1
+ vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a22o_1
XANTENNA__13042__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16160_ clknet_leaf_142_wb_clk_i _01829_ _00389_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\]
+ sky130_fd_sc_hd__dfrtp_1
X_13372_ _07795_ _07797_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__and4b_1
XANTENNA_input86_A wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10584_ team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] net1096 net1053 vssd1 vssd1 vccd1
+ vccd1 _06128_ sky130_fd_sc_hd__and3_1
XFILLER_0_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload19 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15111_ net1139 vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_156_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12323_ net244 net671 vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16091_ clknet_leaf_92_wb_clk_i _01760_ _00320_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12482__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09267__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ net1255 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__inv_2
XANTENNA__08171__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ net245 net673 vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08024__X _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _06604_ _06618_ net554 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__mux2_1
X_12185_ net260 net648 vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11451__S0 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_X net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ net706 _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_79_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16993_ clknet_leaf_131_wb_clk_i _02662_ _01222_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\]
+ sky130_fd_sc_hd__dfrtp_1
X_15944_ clknet_leaf_57_wb_clk_i _01621_ _00171_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__dfrtp_1
X_11067_ net593 net549 vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__and2_1
XANTENNA__12320__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _05588_ _05628_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__or2_1
X_15875_ clknet_leaf_96_wb_clk_i _01552_ _00102_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14826_ net1112 vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__inv_2
XANTENNA__12608__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14757_ net1111 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__inv_2
X_11969_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[2\] team_04_WB.instance_to_wrap.CPU_DAT_O\[2\]
+ net266 vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__mux2_1
XANTENNA__13281__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13708_ net755 _06915_ net271 _07696_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__a31o_1
XANTENNA__08383__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_88_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11831__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14688_ net1213 vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__inv_2
XANTENNA__08346__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13639_ net1001 _03024_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_1
XANTENNA__13033__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16427_ clknet_leaf_30_wb_clk_i _02096_ _00656_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10177__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16358_ clknet_leaf_17_wb_clk_i _02027_ _00587_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[331\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08686__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ net1201 vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14083__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16289_ clknet_leaf_130_wb_clk_i _01958_ _00518_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17261__1321 vssd1 vssd1 vccd1 vccd1 _17261__1321/HI net1321 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_4_11__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09177__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08081__S net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09635__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13887__A2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_97_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09801_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\]
+ net890 vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__mux2_1
Xfanout217 _07277_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__clkbuf_2
Xfanout228 _07438_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_2
XFILLER_0_157_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07993_ _03601_ _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__nand2_1
Xfanout239 _07301_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_52_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ net666 _05342_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12847__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__D net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08515__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09663_ _05270_ _05271_ _05272_ _05273_ net795 net813 vssd1 vssd1 vccd1 vccd1 _05274_
+ sky130_fd_sc_hd__mux4_1
X_08614_ net720 _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _05201_ _05202_ _05203_ _05204_ net794 net814 vssd1 vssd1 vccd1 vccd1 _05205_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14064__A2 net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13272__A0 net95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08545_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__mux2_1
XANTENNA__08279__B1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ net595 _04083_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12286__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__B _06676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13024__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_A _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_X net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10518__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09794__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ _04635_ _04636_ _04637_ _04638_ net836 net748 vssd1 vssd1 vccd1 vccd1 _04639_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11889__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\] vssd1 vssd1
+ vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\] vssd1 vssd1
+ vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[567\] vssd1 vssd1
+ vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_72_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold293 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\] vssd1 vssd1
+ vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09815__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__clkbuf_4
Xfanout762 _03570_ vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__clkbuf_4
Xfanout773 net777 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12838__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _04695_ net263 _03325_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__and3_1
Xfanout784 net790 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
XANTENNA__12302__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout795 net799 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__clkbuf_4
X_12941_ net256 net2286 net321 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_161_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11510__B1 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16010__Q team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__X _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15660_ net1174 vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
X_12872_ _07572_ net338 net388 net2116 vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09550__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ net1226 vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13263__A0 net73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ net704 _05841_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__nor2_1
X_15591_ net1139 vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__inv_2
XANTENNA__13072__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330_ net1386 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
X_14542_ net1263 vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__inv_2
X_11754_ net758 _05544_ net697 _03645_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__a22o_1
XANTENNA__11813__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08166__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_7__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17261_ net1321 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
X_10705_ _06188_ net1057 _05111_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or3b_4
XFILLER_0_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13015__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14473_ net1251 vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ _06217_ _06247_ _06272_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16212_ clknet_leaf_2_wb_clk_i _01881_ _00441_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\]
+ sky130_fd_sc_hd__dfrtp_1
X_13424_ _07739_ _07742_ _07848_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17192_ clknet_leaf_79_wb_clk_i _02804_ _01421_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10636_ _03517_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nor2_8
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output192_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload108 clknet_leaf_114_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload108/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16143_ clknet_leaf_185_wb_clk_i _01812_ _00372_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload119 clknet_leaf_137_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__inv_6
X_13355_ _07778_ _07780_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10567_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[11\]
+ _06116_ net1048 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ net2205 net500 _07597_ net445 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ clknet_leaf_109_wb_clk_i _01743_ _00303_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13286_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ _07714_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__or4_1
X_10498_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\] net1006 _06043_ _06053_
+ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__a22o_1
X_15025_ net1266 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__inv_2
X_12237_ net2329 net504 _07561_ net445 vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a22o_1
XANTENNA__08745__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ net1960 net508 _07525_ net441 vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a22o_1
XANTENNA__13247__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _06241_ _06607_ _06603_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12151__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12829__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16976_ clknet_leaf_192_wb_clk_i _02645_ _01205_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12099_ net2307 net352 _07504_ net443 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a22o_1
X_15927_ clknet_leaf_70_wb_clk_i _01604_ _00154_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_X clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 DAT_I[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14867__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__B1 _05139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15798__17 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__inv_2
X_15858_ clknet_leaf_98_wb_clk_i _01535_ _00085_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13254__A0 net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net1248 vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14078__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11291__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08330_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[762\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__mux2_1
XANTENNA__11804__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09473__A2 _05083_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08261_ net772 _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__or2_2
XANTENNA__13006__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08108__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08141__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__mux2_1
XANTENNA__08804__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12160__C_N net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10240__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12780__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout390_A _07673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout488_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _03583_ _03584_ _03585_ _03586_ net787 net801 vssd1 vssd1 vccd1 vccd1 _03587_
+ sky130_fd_sc_hd__mux4_1
X_09715_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__mux2_1
XANTENNA__12296__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout655_A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14777__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__X _07242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _05253_ _05254_ _05255_ _05256_ net794 net814 vssd1 vssd1 vccd1 vccd1 _05257_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09370__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13245__A0 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09577_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__mux2_1
XANTENNA__12048__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13796__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08528_ _04113_ _04138_ net662 vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__mux2_2
XANTENNA__12599__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08459_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13548__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13548__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ _06798_ _06247_ _06240_ _06789_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08714__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13012__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10421_ net2665 net1006 vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10545__A team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12220__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13140_ _07574_ net382 net297 net2209 vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a22o_1
XANTENNA__11574__A3 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10352_ net282 _05941_ net1057 vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16005__Q team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ net244 net2423 net305 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__mux2_1
X_10283_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] net1056 _05877_
+ _05880_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__a22o_1
XANTENNA__09545__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ net2437 net518 _07464_ net461 vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a22o_1
XANTENNA_input49_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10__f_wb_clk_i_X clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13067__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16830_ clknet_leaf_129_wb_clk_i _02499_ _01059_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08021__Y _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _05251_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_2
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__buf_2
Xfanout592 _04166_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_4
X_16761_ clknet_leaf_154_wb_clk_i _02430_ _00990_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\]
+ sky130_fd_sc_hd__dfrtp_1
X_13973_ _04243_ net262 net598 _03320_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__a31o_1
XANTENNA__12287__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15712_ net1264 vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__inv_2
X_12924_ net212 net2488 net319 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
X_16692_ clknet_leaf_3_wb_clk_i _02361_ _00921_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09280__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13236__A0 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17260__1320 vssd1 vssd1 vccd1 vccd1 _17260__1320/HI net1320 sky130_fd_sc_hd__conb_1
X_15643_ net1179 vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _07553_ net349 net395 net2626 vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a22o_1
XANTENNA_output205_A net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11806_ net689 _06708_ _07288_ net613 vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__o211a_4
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15574_ net1228 vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ _07513_ net345 net398 net1665 vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
XANTENNA__08972__X _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17313_ net1369 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
X_14525_ net1190 vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__inv_2
X_11737_ _06935_ _06955_ _07206_ _07219_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08663__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17244_ net1304 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ net1292 vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08624__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ net559 _06827_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__nor2_1
XANTENNA__13003__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ _07831_ _07832_ _07746_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__inv_2
X_17175_ clknet_leaf_90_wb_clk_i _02787_ _01404_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14387_ net1450 vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12146__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11599_ _06749_ _07087_ net584 vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16126_ clknet_leaf_142_wb_clk_i _01795_ _00355_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_13338_ net1085 team_04_WB.MEM_SIZE_REG_REG\[12\] team_04_WB.MEM_SIZE_REG_REG\[13\]
+ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__or3b_1
XFILLER_0_52_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12762__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_958 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__A1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10605__D net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13766__A team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ clknet_leaf_175_wb_clk_i _01726_ _00286_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_13269_ net98 net2654 net977 vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08718__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12514__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ net1213 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__inv_2
XANTENNA__13711__B2 _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_33 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08813__S1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16959_ clknet_leaf_159_wb_clk_i _02628_ _01188_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\]
+ sky130_fd_sc_hd__dfrtp_1
X_09500_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[11\] team_04_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ net1010 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09190__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11292__Y _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _05038_ _05039_ _05040_ _05041_ net793 net813 vssd1 vssd1 vccd1 vccd1 _05042_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ _04948_ _04972_ net667 vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_47_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11789__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08313_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09293_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__mux2_1
XANTENNA__12450__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 _07692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08244_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\]
+ net878 vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__mux2_1
XANTENNA_33 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08534__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10636__Y _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__A2 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08175_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[508\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[476\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__mux2_1
XANTENNA__10365__A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_X clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12753__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput140 net140 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
Xoutput151 net151 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12505__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput162 net162 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
Xoutput173 net173 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__clkbuf_4
Xoutput184 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput195 net195 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XANTENNA_fanout772_A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1100_X net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net973 _03568_ vssd1 vssd1 vccd1
+ vccd1 _03570_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08776__Y _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__X _06972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout658_X net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10970_ _04329_ _06457_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__C net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_139_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ _07611_ net486 net408 net1639 vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XANTENNA__11930__Y _07396_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12441__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ _07538_ net493 net419 net1881 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ net2487 net1077 vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11522_ _06502_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_156_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12992__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15290_ net1146 vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__inv_2
XANTENNA__12474__B net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ _03428_ _03429_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ net553 _06738_ _06735_ net567 vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08948__A1 _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _05617_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__or2_1
XANTENNA__12744__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14172_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\]
+ _03385_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__and3_1
XANTENNA__11401__C1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ _06871_ _06872_ net566 vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__mux2_1
X_13123_ _07557_ net373 net295 net1899 vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a22o_1
X_10335_ _03498_ net1076 _05926_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09275__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13054_ _07515_ net380 net308 net2022 vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a22o_1
X_10266_ _05569_ _05570_ _05640_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10722__B _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ net226 net680 vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10197_ _05552_ _05553_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__and2b_1
X_16813_ clknet_leaf_42_wb_clk_i _02482_ _01042_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16744_ clknet_leaf_113_wb_clk_i _02413_ _00973_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\]
+ sky130_fd_sc_hd__dfrtp_1
X_13956_ _03807_ net599 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__and2b_1
XANTENNA__09220__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12907_ _07609_ net347 net387 net2085 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__a22o_1
X_13887_ net1604 net1066 net1039 _03267_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a22o_1
X_16675_ clknet_leaf_125_wb_clk_i _02344_ _00904_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10691__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15626_ net1107 vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12838_ _07536_ net346 net395 net2090 vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12769_ _07496_ net326 net396 net2025 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
X_15557_ net1108 vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__inv_2
XANTENNA__10737__X _06226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_168_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_168_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15041__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08731__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508_ net1260 vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__inv_2
XANTENNA__12983__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15488_ net1212 vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__inv_2
XANTENNA__08354__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17227_ net1433 _02837_ _01481_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\]
+ sky130_fd_sc_hd__dfrtp_4
Xinput20 DAT_I[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput31 DAT_I[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ net1276 vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14880__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput64 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09974__A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12735__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput75 wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_1
X_17158_ clknet_leaf_77_wb_clk_i _02770_ _01387_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold804 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\] vssd1 vssd1
+ vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 wbs_dat_i[25] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_1
XFILLER_0_141_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold815 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\] vssd1 vssd1
+ vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10746__A1 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold826 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\] vssd1 vssd1
+ vccd1 vccd1 net2263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 wbs_dat_i[6] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
Xhold837 _02722_ vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ clknet_leaf_41_wb_clk_i _01778_ _00338_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold848 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\] vssd1 vssd1
+ vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14091__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17089_ clknet_leaf_75_wb_clk_i _02724_ _01318_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_09980_ net631 _04839_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold859 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\] vssd1 vssd1
+ vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[47\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XANTENNA__13160__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08798__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ net663 _04441_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ _04400_ _04401_ _04402_ _04403_ net829 net743 vssd1 vssd1 vccd1 vccd1 _04404_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09116__A1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout353_A _07484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08970__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09345_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout520_A _06197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09868__B net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1262_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13023__X _07680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10807__B _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1050_X net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08158_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout987_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[510\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\]
+ net918 vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09095__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10542__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10051_ _03493_ _03728_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nor2_1
XANTENNA__13151__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08012__B net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13853__B net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15785__4 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__inv_2
X_13810_ net753 _06708_ net272 net709 vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__a31o_1
X_14790_ net1106 vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__inv_2
XANTENNA__12102__X _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ _03130_ _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__and2b_1
XFILLER_0_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ net628 _06439_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10673__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ _03058_ _03062_ net1001 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_123_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16460_ clknet_leaf_107_wb_clk_i _02129_ _00689_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__inv_2
XANTENNA__13206__A3 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _07594_ net487 net410 net2137 vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a22o_1
X_15411_ net1246 vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_62_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16391_ clknet_leaf_165_wb_clk_i _02060_ _00620_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12414__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13080__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15342_ net1207 vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12965__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ net699 _06198_ net650 vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__or3b_1
XFILLER_0_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10717__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11505_ _06504_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__and2_1
X_15273_ net1137 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__inv_2
X_12485_ net2520 net430 net489 _07480_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter_state _06170_
+ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__and2_1
XANTENNA_input71_X net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12717__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17012_ clknet_leaf_1_wb_clk_i _02681_ _01241_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\]
+ sky130_fd_sc_hd__dfrtp_1
X_11436_ net636 _04528_ net357 vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11925__B1 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14155_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\]
+ _03529_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11367_ _06848_ _06851_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _07538_ net377 net301 net1600 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a22o_1
X_10318_ net280 _05910_ net1058 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21o_1
X_14086_ net1502 _06118_ net1033 vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__mux2_1
X_11298_ net532 _06573_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13037_ _07498_ net373 net307 net2014 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a22o_1
XANTENNA__13142__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _05685_ _05686_ _05687_ _05763_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1140 net1141 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_4
Xfanout1151 net1153 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_4
Xfanout1162 net1166 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_2
Xfanout1173 net1181 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__buf_4
Xfanout1184 net1186 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_4
Xfanout1195 net1202 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
X_14988_ net1121 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16727_ clknet_leaf_154_wb_clk_i _02396_ _00956_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\]
+ sky130_fd_sc_hd__dfrtp_1
X_13939_ _03057_ _03084_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09969__A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16658_ clknet_leaf_7_wb_clk_i _02327_ _00887_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15609_ net1248 vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12405__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16589_ clknet_leaf_29_wb_clk_i _02258_ _00818_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\]
+ net882 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\]
+ net874 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08012_ _03597_ net905 _03617_ _03620_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold601 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\] vssd1 vssd1
+ vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08812__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold612 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\] vssd1 vssd1
+ vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\] vssd1 vssd1
+ vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07936__B net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[89\] vssd1 vssd1
+ vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\] vssd1 vssd1
+ vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\] vssd1 vssd1
+ vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold667 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\] vssd1 vssd1
+ vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_107_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09963_ _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__nor2_1
Xhold678 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\] vssd1 vssd1
+ vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09209__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_38_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold689 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1006\] vssd1 vssd1
+ vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13133__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13954__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _04519_ _04524_ net722 vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1010_A _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ net639 _04246_ _04302_ _04300_ _04273_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__a32o_1
XANTENNA__09643__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[17\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout470_A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout568_A _05251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ net782 net702 _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a21oi_4
XPHY_EDGE_ROW_108_Left_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout735_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10655__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout902_A net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1265_X net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10407__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_836 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09328_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11604__C1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10958__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_146_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09259_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_519 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_117_Left_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09818__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12270_ net253 net672 vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__and2_1
XANTENNA__08722__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout892_X net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ net753 _06708_ _06686_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13200__Y _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10186__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12580__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _06264_ _06639_ _06640_ net530 vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__o22a_1
XANTENNA__08023__A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _04893_ vssd1
+ vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2_1
XANTENNA__13124__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15960_ clknet_leaf_71_wb_clk_i _01636_ _00189_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11083_ net579 net551 vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__nand2_1
XANTENNA__11135__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__B2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A2 _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12332__B1 _07610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input31_A DAT_I[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08000__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _05564_ _05643_ _05565_ _05563_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__a211o_1
X_14911_ net1265 vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__inv_2
XANTENNA__15852__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15891_ clknet_leaf_99_wb_clk_i _01568_ _00118_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__dfrtp_1
XANTENNA__13075__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14842_ net1146 vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12199__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09187__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11985_ _07398_ _07442_ _07441_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a21o_1
X_14773_ net1200 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09500__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16512_ clknet_leaf_135_wb_clk_i _02181_ _00741_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\]
+ sky130_fd_sc_hd__dfrtp_1
X_13724_ net995 _03112_ _03114_ _07691_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__a22o_1
X_10936_ _06387_ _06390_ _06386_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__o21ba_1
XANTENNA_clkbuf_leaf_185_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_151_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09141__X _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16443_ clknet_leaf_101_wb_clk_i _02112_ _00672_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\]
+ sky130_fd_sc_hd__dfrtp_1
X_13655_ _07103_ net274 _07697_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__o21ai_1
X_10867_ _04528_ _06296_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12606_ _07575_ net493 net414 net1993 vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a22o_1
X_13586_ net992 _02973_ _02976_ net989 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o22a_1
XFILLER_0_143_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11550__C _07037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16374_ clknet_leaf_10_wb_clk_i _02043_ _00603_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ _04974_ _06269_ _06283_ _06285_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15325_ net1149 vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__inv_2
X_12537_ net2241 net259 net421 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15256_ net1205 vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__inv_2
X_12468_ net522 net606 _07469_ net428 net1990 vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a32o_1
XANTENNA__13899__B1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14207_ net1087 _03409_ _03403_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__o21ai_1
X_11419_ net585 _06648_ _06886_ _06643_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_1_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15187_ net1233 vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__inv_2
XANTENNA__12154__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ net2111 net434 _07628_ net523 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12571__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1090
+ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__or2_1
XANTENNA__13115__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09971__B _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ net1464 _06084_ net1033 vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10334__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _04237_ _04238_ _04239_ _04240_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04241_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10885__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08561_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13713__S net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_183_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_183_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_18_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11834__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08807__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_174_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08890__X _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_690 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09044_ net782 _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__nor2_1
XANTENNA__13668__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13020__Y _07679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold420 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\] vssd1 vssd1
+ vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[338\] vssd1 vssd1
+ vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11365__A1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1225_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold442 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\] vssd1 vssd1
+ vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\] vssd1 vssd1
+ vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold464 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\] vssd1 vssd1
+ vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[488\] vssd1 vssd1
+ vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold486 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\] vssd1 vssd1
+ vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
Xhold497 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\] vssd1 vssd1
+ vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net913 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13106__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__B net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout922 net925 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__buf_4
XANTENNA__14132__X net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ net641 _04003_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_74_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout933 net934 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__clkbuf_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__clkbuf_4
Xfanout955 net956 vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__clkbuf_2
Xfanout966 net971 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_4
Xfanout977 net978 vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10325__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__B _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _04586_ _04644_ _05487_ _04585_ _04557_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout852_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1120 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[268\] vssd1 vssd1
+ vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout988 _07704_ vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_4
Xfanout999 _07686_ vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\] vssd1 vssd1
+ vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\] vssd1 vssd1
+ vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ net768 _04432_ _04438_ _04425_ _04426_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__a32oi_4
Xhold1153 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[896\] vssd1 vssd1
+ vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\] vssd1 vssd1
+ vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1175 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\] vssd1 vssd1
+ vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1186 net115 vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ _04366_ _04367_ _04368_ _04369_ net787 net801 vssd1 vssd1 vccd1 vccd1 _04370_
+ sky130_fd_sc_hd__mux4_1
Xhold1197 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\] vssd1 vssd1
+ vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11770_ net613 _07256_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_120_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10819__Y _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10721_ net579 net548 _06209_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_172_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A2 _07317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__A team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_X net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ net1082 team_04_WB.MEM_SIZE_REG_REG\[28\] vssd1 vssd1 vccd1 vccd1 _07866_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08049__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10652_ net1523 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1
+ vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Left_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13371_ _07792_ _07796_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10583_ _06127_ net1542 net1023 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12322_ net2066 net500 _07605_ net447 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a22o_1
X_15110_ net1103 vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16090_ clknet_leaf_44_wb_clk_i _01759_ _00319_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input79_A wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15847__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15041_ net1188 vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12253_ net2181 net504 _07569_ net448 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11204_ net586 _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nand2_1
X_12184_ net2240 net507 _07533_ net437 vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ net464 _06593_ _06623_ net287 vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a22o_2
X_16992_ clknet_leaf_138_wb_clk_i _02661_ _01221_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input34_X net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15943_ clknet_leaf_57_wb_clk_i _01620_ _00170_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__dfrtp_1
X_11066_ _06547_ _06554_ net559 vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__mux2_1
X_10017_ _05592_ _05625_ _05589_ _05590_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15874_ clknet_leaf_86_wb_clk_i _01551_ _00101_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08080__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14825_ net1136 vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11842__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11816__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14756_ net1168 vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__inv_2
X_11968_ _03631_ _05994_ net1059 net756 vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_169_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09312__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ _03018_ _03093_ _03097_ _03096_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__o31a_2
XFILLER_0_156_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08383__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12149__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ net548 net533 net659 vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11899_ net2112 net529 net452 _07369_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14687_ net1248 vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ clknet_leaf_163_wb_clk_i _02095_ _00655_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\]
+ sky130_fd_sc_hd__dfrtp_1
X_13638_ net1000 _03021_ _03028_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__nand3_1
XFILLER_0_132_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10177__B _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16357_ clknet_leaf_169_wb_clk_i _02026_ _00586_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\]
+ sky130_fd_sc_hd__dfrtp_1
X_13569_ _07763_ _07820_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12792__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15308_ net1122 vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16288_ clknet_leaf_136_wb_clk_i _01957_ _00517_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15239_ net1142 vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09635__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09800_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[321\]
+ net893 vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__mux2_1
Xfanout218 _07277_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_1
X_07992_ net1079 net1029 net1025 _03502_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a31o_1
Xfanout229 _07426_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
XANTENNA__10921__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_163_Right_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09731_ _03639_ _03641_ _05337_ _05339_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__a211o_1
XANTENNA__09399__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\]
+ net955 vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08613_ _04220_ _04221_ _04222_ _04223_ net823 net733 vssd1 vssd1 vccd1 vccd1 _04224_
+ sky130_fd_sc_hd__mux4_1
X_09593_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout266_A _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08544_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\]
+ net918 vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08279__A1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12075__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08475_ net595 _04083_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__nand2_1
XANTENNA__11822__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout433_A _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1175_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13024__A1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09323__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14127__X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout600_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11586__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12783__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09027_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[654\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold250 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\] vssd1 vssd1
+ vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold261 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\] vssd1 vssd1
+ vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\] vssd1 vssd1
+ vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\] vssd1 vssd1
+ vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11927__A _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\] vssd1 vssd1
+ vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12522__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14288__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__clkbuf_8
Xfanout741 net742 vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09929_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\]
+ _05539_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout752 _03629_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkbuf_8
Xfanout763 net764 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__clkbuf_8
Xfanout774 net776 vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 net790 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_4
XFILLER_0_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
X_12940_ net258 net2559 net320 vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_161_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_161_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _07571_ net346 net391 net1969 vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a22o_1
XANTENNA__11662__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ net1237 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__inv_2
X_11822_ net2160 net526 net438 _07302_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__a22o_1
XANTENNA__13263__A1 team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15590_ net1103 vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14541_ net1264 vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__inv_2
X_11753_ team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] net270 net268 vssd1 vssd1 vccd1
+ vccd1 _07242_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11813__A2 _06839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _05111_ _06191_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__or2_1
X_17260_ net1320 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_14472_ net1273 vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__inv_2
X_11684_ net575 _06239_ _07172_ net581 vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ clknet_leaf_184_wb_clk_i _01880_ _00440_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\]
+ sky130_fd_sc_hd__dfrtp_1
X_13423_ _07739_ _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__nand2_1
X_10635_ _06159_ _06170_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__or2_2
XFILLER_0_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ clknet_leaf_78_wb_clk_i _02803_ _01420_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09278__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_158_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA__12774__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ _07773_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__nand2_1
X_16142_ clknet_leaf_28_wb_clk_i _01811_ _00371_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06116_ sky130_fd_sc_hd__and3_1
XANTENNA__08182__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10785__C1 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ _07283_ net669 vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__and2_2
X_13285_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[1\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__or2_1
X_16073_ clknet_leaf_120_wb_clk_i _01742_ _00302_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_10497_ _06051_ _06069_ _06070_ net1006 team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15024_ net1164 vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__inv_2
X_12236_ net217 net673 vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ net219 net649 vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__and2_1
X_11118_ _06604_ _06606_ net560 vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__mux2_1
X_16975_ clknet_leaf_189_wb_clk_i _02644_ _01204_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\]
+ sky130_fd_sc_hd__dfrtp_1
X_12098_ net243 net676 vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_30_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15926_ clknet_leaf_70_wb_clk_i _01603_ _00153_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11049_ net581 _06537_ net288 vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o21a_1
Xinput7 DAT_I[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09983__A_N net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15857_ clknet_leaf_96_wb_clk_i _01534_ _00084_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_88 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13263__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ net1225 vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09553__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14739_ net1226 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09977__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _03867_ _03868_ _03869_ _03870_ net788 net809 vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13006__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08108__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16409_ clknet_leaf_178_wb_clk_i _02078_ _00638_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09305__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14094__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10916__A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12765__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12517__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08197__A0 _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11466__B _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[575\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[543\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout383_A _07679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09714_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__mux2_1
XANTENNA__12296__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09645_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[386\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout550_A _05376_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1292_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09576_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__mux2_1
XANTENNA__12048__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12297__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08527_ _04120_ _04126_ _04137_ net716 vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__a22o_2
XFILLER_0_78_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08458_ net727 _04068_ net712 vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08389_ _03994_ _03999_ net770 vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net1085 net1006 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__and2_1
XANTENNA__09098__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12756__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12220__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10545__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09637__A1_N net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10351_ _05530_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12508__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13070_ _07333_ net2597 net303 vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10282_ net281 _05878_ net1056 vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08730__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13181__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ net244 net684 vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_163_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_163_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16021__Q team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 net575 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__buf_2
X_16760_ clknet_leaf_156_wb_clk_i _02429_ _00989_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout582 net584 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12287__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13972_ net148 net1064 vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__and2_1
Xfanout593 _04112_ vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__buf_2
X_15711_ net1262 vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__inv_2
X_12923_ _07246_ net2605 net319 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__mux2_1
XANTENNA__15860__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16691_ clknet_leaf_184_wb_clk_i _02360_ _00920_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13083__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15642_ net1179 vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12854_ _07552_ net344 net394 net1978 vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__a22o_1
X_11805_ net686 _07287_ _07286_ _07285_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__a211o_1
X_15573_ net1215 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__inv_2
X_12785_ _07512_ net341 net398 net1633 vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11798__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17312_ net1368 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_56_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12995__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ net1190 vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11736_ _06816_ _06817_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08905__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ net1405 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
X_14455_ net1291 vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ net289 _06959_ _07155_ net586 vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12747__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13406_ net1085 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 _07832_
+ sky130_fd_sc_hd__and2_1
X_10618_ _06149_ _06150_ _06151_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__or3_1
X_17174_ clknet_leaf_93_wb_clk_i _02786_ _01403_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14386_ net1477 vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__clkbuf_1
X_11598_ net569 _06941_ _07085_ _07086_ _06251_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16125_ clknet_leaf_130_wb_clk_i _01794_ _00354_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_13337_ team_04_WB.MEM_SIZE_REG_REG\[14\] _07761_ _07762_ vssd1 vssd1 vccd1 vccd1
+ _07763_ sky130_fd_sc_hd__a21o_1
X_10549_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[17\]
+ _06104_ net1048 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10773__A2 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16056_ clknet_leaf_153_wb_clk_i _01725_ _00285_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_13268_ net99 team_04_WB.ADDR_START_VAL_REG\[8\] net977 vssd1 vssd1 vccd1 vccd1 _01638_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13172__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ net1265 vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__inv_2
XANTENNA__13711__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_195 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ net221 net649 vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__and2_1
X_13199_ _03548_ _07687_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__and2_1
XFILLER_0_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16958_ clknet_leaf_129_wb_clk_i _02627_ _01187_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09471__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ clknet_leaf_35_wb_clk_i _01586_ _00136_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__dfrtp_1
XANTENNA__14089__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16889_ clknet_leaf_152_wb_clk_i _02558_ _01118_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12398__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13227__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ net718 _04971_ _04960_ _04959_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_47_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08312_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__mux2_1
XANTENNA__11789__B2 _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12986__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12450__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_23 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_34 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10646__A _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12738__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08174_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\]
+ net857 vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12202__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1040_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1138_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput130 net130 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput141 net141 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_101_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout598_A net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 net152 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput163 net163 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
Xoutput174 net174 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput185 net185 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput196 net196 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__buf_2
XANTENNA__12910__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout765_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net973 _03568_ vssd1 vssd1 vccd1
+ vccd1 _03569_ sky130_fd_sc_hd__o21a_1
XANTENNA__12269__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09381__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08568__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__B net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11477__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout932_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\] vssd1 vssd1
+ vccd1 vccd1 _03504_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__mux2_1
XANTENNA__13823__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_52_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09559_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\]
+ net889 vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11940__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15412__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12570_ _07537_ net484 net417 net1799 vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12441__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_156_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ team_04_WB.MEM_SIZE_REG_REG\[6\] _06501_ team_04_WB.MEM_SIZE_REG_REG\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_156_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__Y _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14028__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__C net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12729__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14240_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\] _03426_ net819
+ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__o21ai_1
X_11452_ _06939_ _06940_ net562 vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__mux2_1
Xwire235 _07408_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire257 _07362_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__buf_2
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10403_ _05608_ _05609_ _05616_ net617 vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a31o_1
X_14171_ _03387_ _03388_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08948__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ _06641_ _06714_ net557 vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input61_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ net282 _05925_ _05924_ net1057 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ net700 _07555_ _07666_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__or3_4
XFILLER_0_104_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15855__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_131_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13154__B1 net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13078__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ _07514_ net379 net309 net1732 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10265_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] net1055 _05859_
+ _05864_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a22o_1
XANTENNA__12901__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ net2399 net516 _07455_ net446 vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
XANTENNA__14329__S0 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10196_ _05771_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14103__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ clknet_leaf_119_wb_clk_i _02481_ _01041_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_91_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09291__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout390 _07673_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16743_ clknet_leaf_21_wb_clk_i _02412_ _00972_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\]
+ sky130_fd_sc_hd__dfrtp_1
X_13955_ _03860_ net266 net599 _03311_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkload7_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ _07608_ net350 net386 net2614 vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a22o_1
X_16674_ clknet_leaf_147_wb_clk_i _02343_ _00903_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[647\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12011__A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ _02933_ _03259_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ net1132 vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__inv_2
X_12837_ _07535_ net334 net393 net1769 vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12968__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15556_ net1172 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__inv_2
X_12768_ _07495_ net326 net396 net1812 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14507_ net1260 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__inv_2
X_11719_ _06996_ _07009_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12157__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08731__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ net1273 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
X_12699_ net2143 net404 net329 _07296_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17226_ net1432 _02836_ _01479_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput10 DAT_I[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ net1272 vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 DAT_I[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput32 DAT_I[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput43 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput54 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13777__A team_04_WB.ADDR_START_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12196__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17157_ clknet_leaf_78_wb_clk_i _02769_ _01386_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput65 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14369_ net1510 vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__clkbuf_1
Xhold805 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\] vssd1 vssd1
+ vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xinput76 wbs_dat_i[16] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold816 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\] vssd1 vssd1
+ vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_1
XANTENNA__11943__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput98 wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09466__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_137_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold827 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[489\] vssd1 vssd1
+ vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ clknet_leaf_111_wb_clk_i _01777_ _00337_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11568__Y _07057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08370__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold838 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\] vssd1 vssd1
+ vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_161_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17088_ clknet_leaf_76_wb_clk_i net1702 _01317_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08223__X _03834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold849 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\] vssd1 vssd1
+ vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13145__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08930_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__mux2_1
X_16039_ clknet_leaf_24_wb_clk_i _01708_ _00268_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08247__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09990__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08861_ net719 _04464_ _04470_ _04458_ net661 vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a311oi_2
XANTENNA__08798__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_21 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08792_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[914\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09413_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[551\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08970__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout346_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1088_A team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12959__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15232__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17323__1379 vssd1 vssd1 vccd1 vccd1 _17323__1379/HI net1379 sky130_fd_sc_hd__conb_1
XFILLER_0_59_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09344_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\]
+ net899 vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__mux2_1
XANTENNA__08545__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11226__A3 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12974__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_136_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout513_A net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08117__Y _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1255_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_151_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08157_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\]
+ net923 vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_151_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09376__S net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\]
+ net918 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout882_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13136__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13687__A1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10050_ _05657_ _05658_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14311__A net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14100__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__B2 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ _03123_ _03126_ _03129_ team_04_WB.ADDR_START_VAL_REG\[9\] vssd1 vssd1 vccd1
+ vccd1 _03131_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10952_ net629 _06439_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__nor2_1
XANTENNA__08410__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_175_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13671_ net991 _03025_ _03059_ _03061_ net993 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__o32a_1
XANTENNA__10673__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_167_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10883_ _06370_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_123_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15410_ net1247 vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _07593_ net487 net410 net1656 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a22o_1
X_16390_ clknet_leaf_17_wb_clk_i _02059_ _00619_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[363\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12414__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15341_ net1201 vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ net2332 _07445_ net423 vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11504_ team_04_WB.MEM_SIZE_REG_REG\[9\] _06503_ vssd1 vssd1 vccd1 vccd1 _06993_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15272_ net1118 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__inv_2
X_12484_ _06194_ _07250_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nor2_1
X_17011_ clknet_leaf_181_wb_clk_i _02680_ _01240_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12178__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13597__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ team_04_WB.instance_to_wrap.final_design.uart.receiving _06172_ _07717_ _03418_
+ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11435_ net585 _06923_ _06669_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14154_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or4_2
X_11366_ _04302_ net364 _06270_ _06852_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13127__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ _05910_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__inv_2
X_13105_ _07537_ net374 net299 net1617 vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11297_ _06657_ _06785_ net463 vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__a21o_1
X_14085_ net1480 _06116_ net1033 vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10248_ _05685_ _05686_ _05687_ _05763_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__nor4_1
XANTENNA__11689__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13036_ _07497_ net374 net307 net1839 vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__a22o_1
Xfanout1130 net1131 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__buf_4
Xfanout1141 net1157 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12350__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10179_ _05549_ _05653_ _05786_ net619 vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__a31o_1
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_4
Xfanout1163 net1165 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__buf_4
Xfanout1174 net1181 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_4
Xfanout1185 net1186 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_2
Xfanout1196 net1202 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__buf_2
X_14987_ net1161 vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__inv_2
X_16726_ clknet_leaf_13_wb_clk_i _02395_ _00955_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\]
+ sky130_fd_sc_hd__dfrtp_1
X_13938_ _03088_ net1040 _03301_ net1072 net1676 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_918 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16657_ clknet_leaf_176_wb_clk_i _02326_ _00886_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\]
+ sky130_fd_sc_hd__dfrtp_1
X_13869_ _03200_ _03220_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15608_ net1221 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12405__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16588_ clknet_leaf_110_wb_clk_i _02257_ _00817_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15539_ net1232 vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10967__A2 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09060_ net702 _04669_ _04386_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_127_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09985__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ _03598_ _03608_ _03616_ _03619_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__and4_2
X_17209_ net1415 _02819_ _01445_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08468__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11916__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold602 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\] vssd1 vssd1
+ vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\] vssd1 vssd1
+ vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\] vssd1 vssd1
+ vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\] vssd1 vssd1
+ vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07936__C net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08662__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\] vssd1 vssd1
+ vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13118__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\] vssd1 vssd1
+ vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold668 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\] vssd1 vssd1
+ vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _05572_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold679 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\] vssd1 vssd1
+ vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08913_ _04520_ _04521_ _04522_ _04523_ net828 net743 vssd1 vssd1 vccd1 vccd1 _04524_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13954__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09893_ net594 _04139_ _04166_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout296_A net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08844_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__mux2_1
XANTENNA__10352__B1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12892__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08775_ _03641_ _03644_ _03640_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_4
XANTENNA_fanout463_A _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12644__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10655__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout251_X net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_A _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout728_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10407__A1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_153_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout516_X net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1258_X net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09258_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\]
+ net924 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08209_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[29\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12525__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09189_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1003\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__mux2_1
XANTENNA__10834__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11907__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11220_ net753 _06686_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13109__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ net644 _03891_ net544 vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10102_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nand2_1
X_11082_ net541 _06570_ _05476_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__a21oi_1
X_10033_ _05564_ _05643_ _05565_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__a21o_1
XANTENNA__12332__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ net1239 vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__inv_2
XANTENNA__15137__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15890_ clknet_leaf_124_wb_clk_i _01567_ _00117_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12883__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A DAT_I[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ net1244 vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14976__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14772_ net1208 vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__inv_2
XANTENNA__09187__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[0\] team_04_WB.instance_to_wrap.CPU_DAT_O\[0\]
+ net266 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__mux2_1
XANTENNA__12635__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16511_ clknet_leaf_160_wb_clk_i _02180_ _00740_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\]
+ sky130_fd_sc_hd__dfrtp_1
X_13723_ _03499_ _05941_ net1102 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
X_10935_ _06392_ _06396_ _06422_ _06390_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ clknet_leaf_39_wb_clk_i _02111_ _00671_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _03043_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08185__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10866_ _06346_ _06350_ _06354_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12399__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _07574_ net492 net415 net2218 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ clknet_leaf_34_wb_clk_i _02042_ _00602_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\]
+ sky130_fd_sc_hd__dfrtp_1
X_13585_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] _05920_ net1100
+ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ _06269_ _06283_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nor3_2
XFILLER_0_54_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15324_ net1148 vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__inv_2
X_12536_ net2495 net244 net423 vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15255_ net1230 vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__inv_2
X_12467_ net525 net607 _07468_ net431 net1703 vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14206_ _03409_ _03410_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_144_Right_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _04814_ _06248_ net362 _04813_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__a221o_1
X_15186_ net1246 vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__inv_2
X_12398_ net653 net609 net219 vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14137_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] _03359_
+ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] vssd1 vssd1 vccd1
+ vccd1 _03360_ sky130_fd_sc_hd__or3b_1
X_11349_ _06279_ _06824_ _06835_ _06837_ net286 vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17322__1378 vssd1 vssd1 vccd1 vccd1 _17322__1378/HI net1378 sky130_fd_sc_hd__conb_1
X_14068_ net1484 _06082_ net1034 vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__mux2_1
XANTENNA__13266__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _07654_ net472 net313 net2349 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_33_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12874__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08560_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\]
+ net851 vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
XANTENNA__12626__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10637__A1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16709_ clknet_leaf_4_wb_clk_i _02378_ _00938_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\]
+ sky130_fd_sc_hd__dfrtp_1
X_08491_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\]
+ net911 vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13051__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__C1 _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _04705_ _04711_ _04722_ net767 vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__a22o_2
XFILLER_0_174_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_152_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_152_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13949__B net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08823__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09043_ _04650_ _04651_ _04652_ _04653_ net789 net801 vssd1 vssd1 vccd1 vccd1 _04654_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout211_A _07246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout309_A _07680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[122\] vssd1 vssd1
+ vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold421 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\] vssd1 vssd1
+ vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\] vssd1 vssd1
+ vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[637\] vssd1 vssd1
+ vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold454 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\] vssd1 vssd1
+ vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold465 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\] vssd1 vssd1
+ vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1120_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[105\] vssd1 vssd1
+ vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold487 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\] vssd1 vssd1
+ vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09654__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold498 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\] vssd1 vssd1
+ vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 net902 vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_4
X_09945_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__nand2b_1
Xfanout912 net913 vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15953__Q team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 net925 vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout580_A _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout934 net941 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 net950 vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_A net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12314__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net962 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ net634 _04698_ _04754_ _05486_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a31o_1
XANTENNA__08613__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
Xfanout978 _07708_ vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12865__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1110 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\] vssd1 vssd1
+ vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout989 net991 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_2
Xhold1121 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\] vssd1 vssd1
+ vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 net110 vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ net781 _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__or2_1
Xhold1143 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\] vssd1 vssd1
+ vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 team_04_WB.instance_to_wrap.final_design.uart.working_data\[7\] vssd1 vssd1
+ vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1165 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\] vssd1 vssd1
+ vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[275\] vssd1 vssd1
+ vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1187 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[320\] vssd1 vssd1
+ vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[18\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1198 team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\] vssd1 vssd1 vccd1
+ vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12617__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08689_ _04274_ _04299_ net662 vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_2
XFILLER_0_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ net625 net551 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10651_ net1548 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1
+ vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _07790_ _07791_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__and2b_1
X_10582_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[6\]
+ _06126_ net1050 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ net245 net669 vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__and2_2
XFILLER_0_146_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12482__C net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ net1213 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12252_ net260 net673 vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__and2_1
XANTENNA__12553__A1 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net574 _06691_ _06532_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a21oi_1
X_12183_ net246 net647 vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__and2_1
XANTENNA__08852__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11134_ net581 _06608_ _06622_ _06599_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__o211a_1
X_16991_ clknet_leaf_159_wb_clk_i _02660_ _01220_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15863__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07980__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13086__S net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11395__A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15942_ clknet_leaf_57_wb_clk_i _01619_ _00169_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__dfrtp_1
X_11065_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__inv_2
X_10016_ _05590_ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and2_1
X_15873_ clknet_leaf_87_wb_clk_i _01550_ _00100_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08080__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14058__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12003__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14824_ net1124 vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13805__A1 team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14755_ net1182 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__inv_2
XANTENNA__11816__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ net2366 net528 net456 _07427_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a22o_1
XANTENNA__10739__A _06227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ _03005_ _03095_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__nand2_1
XANTENNA__11292__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10918_ net625 _06405_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__xnor2_1
X_14686_ net1214 vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11898_ net655 _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__and2_1
X_16425_ clknet_leaf_102_wb_clk_i _02094_ _00654_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\]
+ sky130_fd_sc_hd__dfrtp_1
X_13637_ net991 _03027_ net993 vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13033__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ _06336_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ clknet_leaf_167_wb_clk_i _02025_ _00585_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\]
+ sky130_fd_sc_hd__dfrtp_1
X_13568_ _07151_ net273 _07697_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13769__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10252__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15307_ net1122 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12519_ _07516_ net492 net427 net1729 vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16287_ clknet_leaf_161_wb_clk_i _01956_ _00516_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[260\]
+ sky130_fd_sc_hd__dfrtp_1
X_13499_ net1092 _02889_ net1043 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15238_ net1104 vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__inv_2
XFILLER_0_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12544__A1 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11857__X _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09982__B net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15169_ net1130 vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout219 net220 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_2
X_07991_ net1078 net1030 net1026 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__o31a_1
X_09730_ _03643_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_52_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09399__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10307__B1 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12847__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14049__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08612_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[276\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
X_09592_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08818__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08543_ net779 _04153_ _04148_ net761 vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__o211a_1
X_15812__31 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__inv_2
XFILLER_0_49_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08474_ net595 _04083_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13024__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1070_A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout426_A net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09649__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09323__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08987__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout795_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12535__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13732__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold240 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\] vssd1 vssd1
+ vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12803__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\] vssd1 vssd1
+ vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_X net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_148_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold262 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\] vssd1 vssd1
+ vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09384__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold273 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\] vssd1 vssd1
+ vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold284 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[631\] vssd1 vssd1
+ vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08141__X _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold295 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\] vssd1 vssd1
+ vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout962_A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net723 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout731 net732 vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _05538_ vssd1
+ vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and2_1
Xfanout742 net750 vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__clkbuf_8
Xfanout753 net755 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12104__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12838__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout764 _03570_ vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_4
Xfanout775 net776 vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
Xfanout786 net790 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_8
X_09859_ _04784_ _05456_ _05468_ _03621_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__a22o_2
Xfanout797 net798 vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_161_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _07570_ net336 net389 net1868 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a22o_1
XANTENNA__11662__B _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ net652 net239 vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and2_1
X_14540_ net1286 vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__inv_2
XANTENNA__11274__A1 _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] _07236_ _07240_ _07239_ vssd1
+ vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__a31o_1
XANTENNA__12471__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16019__Q team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ _05111_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__nor2_2
X_14471_ net1250 vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__inv_2
XANTENNA__13015__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11683_ net573 _06224_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nor2_1
X_17321__1377 vssd1 vssd1 vccd1 vccd1 _17321__1377/HI net1377 sky130_fd_sc_hd__conb_1
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16210_ clknet_leaf_7_wb_clk_i _01879_ _00439_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[183\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13422_ _07736_ _07847_ _07738_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input91_A wbs_dat_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09559__S net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17190_ clknet_leaf_78_wb_clk_i _02802_ _01419_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ _06170_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15858__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16141_ clknet_leaf_41_wb_clk_i _01810_ _00370_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\]
+ sky130_fd_sc_hd__dfrtp_1
X_13353_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] team_04_WB.MEM_SIZE_REG_REG\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ _06115_ net1574 net1020 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ net2141 net500 _07596_ net445 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ clknet_leaf_110_wb_clk_i _01741_ _00301_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[3\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[8\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__or4_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10496_ _06036_ _06044_ _06049_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__or3_1
XFILLER_0_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output178_A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15023_ net1140 vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__inv_2
X_12235_ net2270 net504 _07560_ net441 vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ net1974 net509 _07524_ net450 vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
XANTENNA__07953__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ net537 _06235_ _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16974_ clknet_leaf_42_wb_clk_i _02643_ _01203_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\]
+ sky130_fd_sc_hd__dfrtp_1
X_12097_ net2540 net355 _07503_ net452 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
XANTENNA__12829__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ clknet_leaf_70_wb_clk_i _01602_ _00152_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfrtp_2
X_11048_ _06536_ _06532_ _06530_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__or3b_1
Xinput8 DAT_I[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_15856_ clknet_leaf_96_wb_clk_i _01533_ _00083_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_14807_ net1228 vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__inv_2
X_12999_ _07648_ net469 net310 net2262 vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14738_ net1237 vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__inv_2
XANTENNA__12462__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14669_ net1210 vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09469__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16408_ clknet_leaf_150_wb_clk_i _02077_ _00637_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15060__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08190_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
XANTENNA__09305__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08373__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16339_ clknet_leaf_182_wb_clk_i _02008_ _00568_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12690__Y _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_144_Left_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08197__A1 _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09057__X _04668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__B net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07974_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13470__A1_N net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09713_ net776 _05317_ net764 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o21ai_1
XANTENNA__13962__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_A net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_153_Left_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08526_ _04131_ _04136_ net727 vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10098__B _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout710_A _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__Y _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08457_ _04064_ _04065_ _04066_ _04067_ net825 net734 vssd1 vssd1 vccd1 vccd1 _04068_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout808_A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08388_ _03995_ _03996_ _03997_ _03998_ net783 net800 vssd1 vssd1 vccd1 vccd1 _03999_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13953__B1 _03310_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_162_Left_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10545__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10350_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05529_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_115_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12508__A1 _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09009_ net1008 net1007 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\]
+ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_167_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10281_ _05878_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__inv_2
XANTENNA__11938__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12533__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10842__A _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12020_ net2481 net516 _07463_ net447 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__a22o_1
XANTENNA__09480__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_163_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07935__A1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07935__B2 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout550 _05376_ vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_81_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14130__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout561 _05309_ vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11944__Y _07408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout572 net575 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
X_13971_ _04299_ net262 net598 _03319_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__a31o_1
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
Xfanout594 _04112_ vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_171_Left_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15710_ net1281 vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__inv_2
XANTENNA__11673__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _07249_ _07666_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__or2_4
X_16690_ clknet_leaf_10_wb_clk_i _02359_ _00919_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[663\]
+ sky130_fd_sc_hd__dfrtp_1
X_15641_ net1177 vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__inv_2
XANTENNA__09143__A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _07551_ net344 net394 net1801 vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11804_ team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] net270 net268 vssd1 vssd1 vccd1
+ vccd1 _07287_ sky130_fd_sc_hd__a21o_1
X_15572_ net1236 vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__inv_2
X_12784_ _07511_ net342 net398 net2410 vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a22o_1
X_17311_ net1367 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
X_14523_ net1186 vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__inv_2
XFILLER_0_173_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12995__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11735_ _07151_ _07152_ _07222_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08663__A2 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17242_ net1303 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input94_X net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14454_ net1291 vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11666_ _06535_ _06967_ _06252_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ net1084 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 _07831_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10207__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13944__B1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10617_ _06140_ _06146_ _06153_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and3_1
X_17173_ clknet_leaf_93_wb_clk_i _02785_ _01402_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09612__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14385_ net1493 vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ net565 _07028_ net578 vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ clknet_leaf_128_wb_clk_i _01793_ _00353_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\]
+ sky130_fd_sc_hd__dfrtp_1
X_13336_ _07756_ _07760_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10548_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net1094 net1052 vssd1 vssd1 vccd1
+ vccd1 _06104_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16055_ clknet_leaf_166_wb_clk_i _01724_ _00284_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_13267_ net100 net2661 net977 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__mux2_1
X_10479_ _06013_ _06047_ _06050_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or3b_1
XFILLER_0_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15006_ net1218 vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__inv_2
X_12218_ net2422 net509 _07550_ net456 vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a22o_1
XANTENNA__09318__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _07688_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__nand2_1
XANTENNA__07926__A1 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ net252 net2548 net512 vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09752__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14121__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16957_ clknet_leaf_131_wb_clk_i _02626_ _01186_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13274__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1026 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15055__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12683__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ clknet_leaf_11_wb_clk_i _01585_ _00135_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08368__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16888_ clknet_leaf_150_wb_clk_i _02557_ _01117_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12398__B net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15839_ clknet_leaf_90_wb_clk_i _01516_ _00066_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09988__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _04965_ _04970_ net730 vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08311_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[137\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_126_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12450__A3 _07455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_13 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09199__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08242_ _03849_ _03850_ _03851_ _03852_ net831 net747 vssd1 vssd1 vccd1 vccd1 _03853_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_24 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08173_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\]
+ net856 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_95_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11410__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__B2 _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 net120 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__clkbuf_4
XANTENNA__14134__A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput131 net131 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1033_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput142 net142 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput153 net153 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput164 net164 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
Xoutput175 net175 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout493_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput186 net186 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput197 net197 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__buf_2
X_17320__1376 vssd1 vssd1 vccd1 vccd1 _17320__1376/HI net1376 sky130_fd_sc_hd__conb_1
XANTENNA__14112__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[19\] net1009
+ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10601__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\] vssd1 vssd1
+ vccd1 vccd1 _03503_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_165_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_168_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1190_X net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1288_X net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09898__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09558_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[37\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__mux2_1
XANTENNA__12977__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ net720 _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12528__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__mux2_1
XANTENNA__10837__A _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11520_ net708 _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14028__B team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire225 _07414_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__clkbuf_2
X_11451_ net634 _04724_ net630 net632 net552 net540 vssd1 vssd1 vccd1 vccd1 _06940_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10402_ net2643 net1058 _05985_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a21bo_1
X_14170_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _03385_
+ _03381_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11401__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11382_ _06715_ _06870_ net557 vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__mux2_1
X_13121_ _07553_ net382 net301 net1792 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\] _05531_ vssd1
+ vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10572__A team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input54_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _07513_ net379 net308 net1650 vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__a22o_1
X_10264_ _05642_ net620 _05860_ _05863_ net280 vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__a311o_1
XANTENNA__08042__A team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09453__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14979__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ net227 net681 vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__and2_1
XANTENNA__08030__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14329__S1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__nand2b_1
XANTENNA__14103__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16811_ clknet_leaf_15_wb_clk_i _02480_ _01040_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15871__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout391 _07673_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_2
XANTENNA__11468__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16742_ clknet_leaf_22_wb_clk_i _02411_ _00971_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\]
+ sky130_fd_sc_hd__dfrtp_1
X_13954_ net157 net1070 vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08188__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ _07607_ net338 net385 net1670 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a22o_1
XANTENNA_output210_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16673_ clknet_leaf_135_wb_clk_i _02342_ _00902_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\]
+ sky130_fd_sc_hd__dfrtp_1
X_13885_ net1039 _03262_ _03266_ net1068 net1641 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a32o_1
XANTENNA__12011__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12836_ _07534_ net339 net393 net1671 vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a22o_1
X_15624_ net1116 vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__inv_2
XANTENNA__12417__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12968__A1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15555_ net1172 vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13090__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ _07494_ net329 net396 net1830 vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10747__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14506_ net1259 vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__inv_2
X_11718_ _06932_ _06934_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11640__A1 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15486_ net1236 vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12698_ net1903 net404 net327 _07290_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17225_ net1431 _02835_ _01477_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\]
+ sky130_fd_sc_hd__dfrtp_2
X_14437_ net1276 vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ _07011_ _07024_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__xor2_1
Xinput11 DAT_I[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput22 DAT_I[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XANTENNA__09747__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 DAT_I[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
X_17156_ clknet_leaf_73_wb_clk_i _02768_ _01385_ vssd1 vssd1 vccd1 vccd1 team_04_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput55 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08651__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14368_ net1472 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__clkbuf_1
Xinput66 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_1
Xinput77 wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_1
Xhold806 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\] vssd1 vssd1
+ vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13269__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold817 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\] vssd1 vssd1
+ vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ clknet_leaf_23_wb_clk_i _01776_ _00336_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_13319_ team_04_WB.MEM_SIZE_REG_REG\[21\] _07744_ vssd1 vssd1 vccd1 vccd1 _07745_
+ sky130_fd_sc_hd__nand2_1
Xinput88 wbs_dat_i[27] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold828 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\] vssd1 vssd1
+ vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 wbs_dat_i[8] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_2
X_17087_ clknet_leaf_76_wb_clk_i net2274 _01316_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold839 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\] vssd1 vssd1
+ vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
X_14299_ net2037 _03463_ _03465_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09349__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16038_ clknet_leaf_19_wb_clk_i _01707_ _00267_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08247__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__X _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_177_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_177_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08860_ net719 _04464_ _04470_ _04458_ vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__a31o_1
XANTENNA__09482__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_106_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08791_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1010\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12656__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09412_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13081__A0 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout241_A _07295_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_158_Right_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08183__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout339_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09274_ _04881_ _04882_ _04883_ _04884_ net786 net806 vssd1 vssd1 vccd1 vccd1 _04885_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08225_ net752 _03835_ _03725_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__a21o_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1150_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout506_A _07556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ net780 _03766_ net763 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_151_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08087_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\]
+ net918 vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout875_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11698__A1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux2_1
XANTENNA__13990__X _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12647__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10951_ net629 _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13670_ _07795_ _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__nand2_1
XANTENNA__10673__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10882_ _04668_ _06369_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12621_ _07592_ net483 net409 net1749 vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a22o_1
XANTENNA__13072__A0 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15340_ net1129 vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__inv_2
X_12552_ net2468 _07438_ net422 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ net708 _06991_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15271_ net1142 vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12483_ net2379 net430 _07654_ net524 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a22o_1
X_17010_ clknet_leaf_9_wb_clk_i _02679_ _01239_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\]
+ sky130_fd_sc_hd__dfrtp_1
X_14222_ net2652 _06172_ _03418_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a21o_1
XANTENNA__12178__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11434_ _06822_ _06922_ net572 vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__mux2_2
XANTENNA__15866__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11386__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11398__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03372_
+ _03534_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11365_ _04273_ _04301_ net357 _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__o31a_1
XFILLER_0_10_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_13104_ _07536_ net382 net301 net1909 vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a22o_1
X_10316_ _05533_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14084_ net1475 _06114_ net1032 vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__mux2_1
X_11296_ _06350_ _06470_ _06474_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__or3_1
XANTENNA__09426__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13678__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13035_ _07496_ net367 net306 net1706 vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a22o_1
X_10247_ _05643_ _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__xor2_1
XANTENNA__14502__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1120 net1123 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12350__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1131 net1158 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__buf_2
Xfanout1142 net1144 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__buf_4
X_10178_ _05549_ _05653_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a21oi_1
Xfanout1153 net1156 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__buf_4
XANTENNA__14221__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1165 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__buf_2
Xfanout1175 net1181 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__buf_4
Xfanout1186 net1187 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
Xfanout1197 net1202 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
XANTENNA__12638__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ net1106 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16725_ clknet_leaf_12_wb_clk_i _02394_ _00954_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[698\]
+ sky130_fd_sc_hd__dfrtp_1
X_13937_ _03045_ _03086_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nand2_1
XANTENNA__10113__A1 _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13868_ _03250_ _03253_ net1782 net1066 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11861__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16656_ clknet_leaf_190_wb_clk_i _02325_ _00885_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ net1231 vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__inv_2
XANTENNA__13063__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ net230 net2402 net324 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13799_ team_04_WB.ADDR_START_VAL_REG\[16\] _03189_ vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__and2_1
X_16587_ clknet_leaf_16_wb_clk_i _02256_ _00816_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12810__A0 _07374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11074__C1 _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__A1 _06204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15538_ net1247 vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11613__B2 _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13788__A team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15469_ net1143 vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08010_ _03618_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__nor2_4
X_17208_ net1414 _02818_ _01443_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08468__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold603 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[49\] vssd1 vssd1
+ vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_17139_ clknet_leaf_81_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[4\]
+ _01368_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_142_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold614 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\] vssd1 vssd1
+ vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\] vssd1 vssd1
+ vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\] vssd1 vssd1
+ vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold647 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\] vssd1 vssd1
+ vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[335\] vssd1 vssd1
+ vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap366 _04978_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_1
X_09961_ _04440_ _04441_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__nand2_1
Xhold669 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\] vssd1 vssd1
+ vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08912_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[688\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[656\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15508__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _04142_ _04193_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__nor2_1
XANTENNA__12877__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08843_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\]
+ net903 vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__mux2_1
XANTENNA__10352__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08774_ net765 _04377_ _04383_ _04371_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__a31o_2
XANTENNA__12629__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13970__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13841__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11771__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1198_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10655__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13054__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout623_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__mux2_1
XANTENNA__12801__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11604__A1 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09257_ _04814_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12806__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08208_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__mux2_1
XANTENNA__09387__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08291__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09188_ net727 _04798_ net712 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_161_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08139_ _03746_ _03747_ _03748_ _03749_ net831 net747 vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_79_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12580__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ net643 net550 net530 vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _03499_ _04839_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__nand2_1
XANTENNA__08023__C net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ net625 net547 _06569_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__a21o_1
XANTENNA__12868__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12332__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ net639 _04219_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__o21a_1
XANTENNA__11665__B _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ net1225 vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input17_A DAT_I[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ net1226 vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__inv_2
X_11983_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] net759 _03631_
+ _07440_ net696 vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08839__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ net1093 _03112_ net1045 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__o2bb2a_1
X_16510_ clknet_leaf_114_wb_clk_i _02179_ _00739_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ _06392_ _06396_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ team_04_WB.ADDR_START_VAL_REG\[4\] _03042_ vssd1 vssd1 vccd1 vccd1 _03044_
+ sky130_fd_sc_hd__nor2_1
X_16441_ clknet_leaf_178_wb_clk_i _02110_ _00670_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[414\]
+ sky130_fd_sc_hd__dfrtp_1
X_10865_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13596__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12399__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12604_ _07573_ net493 net415 net2082 vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13596__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16372_ clknet_leaf_2_wb_clk_i _02041_ _00601_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\]
+ sky130_fd_sc_hd__dfrtp_1
X_13584_ net998 _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_782 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10796_ _05030_ _05084_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ net1112 vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ net2298 net245 net421 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15254_ net1221 vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__inv_2
X_12466_ net525 net611 _07467_ net431 net1722 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ net1088 _03406_ _03403_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11417_ net633 net590 net358 vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__nor3_1
X_15185_ net1271 vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__inv_2
X_12397_ net2125 net434 _07627_ net523 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a22o_1
XANTENNA__08775__A1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03356_
+ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__or3_1
XANTENNA__12571__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ _04086_ net362 _06257_ _04085_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14067_ net1483 _06080_ net1032 vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__mux2_1
XANTENNA__12859__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _06765_ _06767_ net558 vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08501__Y _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _07653_ net472 net312 net2019 vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a22o_1
XANTENNA__08527__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire257_A _07362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09760__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ net1241 vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__inv_2
XANTENNA__10759__X _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13282__S _05525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16708_ clknet_leaf_169_wb_clk_i _02377_ _00937_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11834__A1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08490_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_56 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16639_ clknet_leaf_157_wb_clk_i _02308_ _00868_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[612\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13036__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09996__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _04716_ _04721_ net774 vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09042_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09000__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_192_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_192_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold400 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\] vssd1 vssd1
+ vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\] vssd1 vssd1
+ vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 net107 vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12562__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\] vssd1 vssd1
+ vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold444 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\] vssd1 vssd1
+ vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_121_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold455 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\] vssd1 vssd1
+ vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\] vssd1 vssd1
+ vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\] vssd1 vssd1
+ vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13457__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09944_ net642 net660 vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__nand2_1
Xhold488 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\] vssd1 vssd1
+ vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout902 net903 vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__buf_4
XANTENNA__12361__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold499 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[225\] vssd1 vssd1
+ vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net926 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__clkbuf_2
Xfanout924 net925 vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net937 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12314__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_A DAT_I[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _04723_ _04753_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__nor2_1
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10325__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1100 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\] vssd1 vssd1
+ vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout968 net971 vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08613__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net981 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__clkbuf_4
Xhold1111 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\] vssd1 vssd1
+ vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\] vssd1 vssd1
+ vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ _04433_ _04434_ _04435_ _04436_ net798 net803 vssd1 vssd1 vccd1 vccd1 _04437_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1133 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\] vssd1 vssd1
+ vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1144 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\] vssd1 vssd1
+ vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\] vssd1 vssd1
+ vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13275__A0 net80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1166 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\] vssd1 vssd1
+ vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08757_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[82\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__mux2_1
Xhold1177 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\] vssd1 vssd1
+ vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\] vssd1 vssd1
+ vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1199 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\] vssd1 vssd1
+ vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11825__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08688_ _04281_ _04287_ _04298_ net716 vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__a22o_4
XANTENNA__08286__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15701__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07978__X _03589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_172_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ net1571 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1
+ vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a22o_1
XANTENNA__08049__A3 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10581_ team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] net1096 net1054 vssd1 vssd1 vccd1
+ vccd1 _06126_ sky130_fd_sc_hd__and3_1
XANTENNA__12536__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10845__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ net2147 net500 _07604_ net447 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ net2395 net503 _07568_ net437 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11202_ net557 _06531_ net356 _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ net2035 net507 _07532_ net436 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a22o_1
XANTENNA__08852__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _06208_ _06621_ _06611_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a21oi_1
X_16990_ clknet_leaf_115_wb_clk_i _02659_ _01219_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\]
+ sky130_fd_sc_hd__dfrtp_1
X_15941_ clknet_leaf_57_wb_clk_i _01618_ _00168_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__dfrtp_1
X_11064_ _06550_ _06552_ net536 vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__mux2_1
XANTENNA__11395__B _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A0 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _05592_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__or2_1
X_15872_ clknet_leaf_87_wb_clk_i _01549_ _00099_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_48_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13266__A0 net70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14823_ net1142 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11816__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11816__B2 _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11966_ net654 net230 vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__and2_1
X_14754_ net1255 vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__inv_2
XANTENNA__10739__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13705_ _03005_ _03015_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_156_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ net625 _06405_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__or2_1
XANTENNA__13018__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685_ net1154 vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11897_ net690 _06899_ _07367_ net614 vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__o211a_2
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13636_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05976_ net1101
+ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
X_16424_ clknet_leaf_112_wb_clk_i _02093_ _00653_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\]
+ sky130_fd_sc_hd__dfrtp_1
X_10848_ net596 _06335_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08924__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ team_04_WB.ADDR_START_VAL_REG\[15\] _02955_ vssd1 vssd1 vccd1 vccd1 _02958_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__08445__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16355_ clknet_leaf_117_wb_clk_i _02024_ _00584_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12241__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10779_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15306_ net1106 vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__inv_2
X_12518_ _07515_ net489 net426 net1972 vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16286_ clknet_leaf_158_wb_clk_i _01955_ _00515_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\]
+ sky130_fd_sc_hd__dfrtp_1
X_13498_ _07858_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15237_ net1110 vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__inv_2
X_12449_ net2581 net429 _07645_ net521 vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15168_ net1211 vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__inv_2
X_14119_ team_04_WB.MEM_SIZE_REG_REG\[18\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[18\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_35_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07990_ _03511_ net1078 net1030 net1026 vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__or4_1
X_15099_ net1113 vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17276__1335 vssd1 vssd1 vccd1 vccd1 _17276__1335/HI net1335 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_52_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14897__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09490__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[372\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08542_ _04149_ _04150_ _04151_ _04152_ net785 net801 vssd1 vssd1 vccd1 vccd1 _04153_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10649__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13009__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ net661 _04081_ _04082_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout321_A _07675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08987__A1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12783__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[526\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1230_A net1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\] vssd1 vssd1
+ vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 net165 vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 net111 vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout690_A net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\] vssd1 vssd1
+ vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold274 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\] vssd1 vssd1
+ vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold285 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[718\] vssd1 vssd1
+ vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold296 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\] vssd1 vssd1
+ vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout710 _07696_ vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__clkbuf_4
Xfanout721 net723 vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__clkbuf_4
Xfanout732 _03667_ vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13982__Y _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09927_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\]
+ _05537_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_165_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13496__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
Xfanout754 net755 vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout955_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net769 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__clkbuf_8
Xfanout776 net777 vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__buf_4
Xfanout787 net788 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_8
X_09858_ _04784_ _05456_ _05468_ _03621_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__a22oi_4
Xfanout798 net799 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09253__X _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__mux2_1
X_11820_ net693 _07182_ _07300_ net615 vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__a211oi_4
XANTENNA__12120__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11751_ _04670_ _05443_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout910_X net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12471__A1 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10702_ net700 _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__or2_2
XANTENNA__10482__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14470_ net1250 vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__inv_2
X_11682_ net581 _07016_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13421_ net1083 team_04_WB.MEM_SIZE_REG_REG\[23\] vssd1 vssd1 vccd1 vccd1 _07847_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10633_ _06160_ _06161_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__or3_2
XFILLER_0_147_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__A team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16140_ clknet_leaf_111_wb_clk_i _01809_ _00369_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_13352_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] team_04_WB.MEM_SIZE_REG_REG\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__nand2_1
XANTENNA__12774__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13971__A1 _04299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input84_A wbs_dat_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[12\]
+ _06114_ net1047 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12303_ net217 net669 vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__and2_1
XANTENNA__11958__X _07420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16071_ clknet_leaf_24_wb_clk_i _01740_ _00300_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_13283_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__or4bb_1
XTAP_TAPCELL_ROW_20_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10495_ _06044_ _06049_ _06036_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_20_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09575__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15022_ net1195 vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12234_ net219 net674 vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__and2_1
XANTENNA__15874__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10514__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ net215 net649 vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08051__Y _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11116_ net537 _06231_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__nor2_1
X_16973_ clknet_leaf_42_wb_clk_i _02642_ _01202_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\]
+ sky130_fd_sc_hd__dfrtp_1
X_12096_ net255 net679 vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15924_ clknet_leaf_70_wb_clk_i _01601_ _00151_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11047_ _06531_ _06534_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__or2_1
XANTENNA__14510__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 DAT_I[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
XANTENNA__13239__A0 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15855_ clknet_leaf_98_wb_clk_i _01532_ _00082_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_14806_ net1221 vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__inv_2
X_12998_ _07647_ net469 net310 net2283 vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ net1267 vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__inv_2
X_11949_ _07398_ _07411_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_116_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_156_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08654__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14668_ net1128 vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__inv_2
XANTENNA__13006__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16407_ clknet_leaf_167_wb_clk_i _02076_ _00636_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08418__A0 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] net1045 _03006_
+ net1098 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12214__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ net1185 vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12765__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16338_ clknet_leaf_10_wb_clk_i _02007_ _00567_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\]
+ sky130_fd_sc_hd__dfrtp_1
X_16269_ clknet_leaf_41_wb_clk_i _01938_ _00498_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_164_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13714__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12517__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13714__B2 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12205__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07973_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[671\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09712_ net781 _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__nor2_1
XANTENNA__12150__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__mux2_1
XANTENNA__11763__B net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_155_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout271_A _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09574_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[613\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08525_ _04132_ _04133_ _04134_ _04135_ net824 net741 vssd1 vssd1 vccd1 vccd1 _04136_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1180_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1278_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08456_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08564__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__X _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08387_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\]
+ net910 vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout324_X net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12756__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12814__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09395__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12508__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ _03504_ net1008 net1007 _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_167_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _05535_ vssd1
+ vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11938__B net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13181__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09480__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net542 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11954__A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14130__B2 team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 net563 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08739__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ net149 net1064 vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__and2_1
XANTENNA__12141__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout573 net574 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_2
Xfanout584 _05140_ vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_2
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_2
X_12921_ _07623_ net349 net387 net2633 vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ net1177 vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__inv_2
X_12852_ _07550_ net345 net394 net1819 vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11803_ net758 _05824_ net697 _04004_ net693 vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__a221o_1
X_12783_ _07510_ net342 net398 net2062 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__a22o_1
X_15571_ net1244 vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17310_ net1366 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
X_14522_ net1186 vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__inv_2
X_11734_ _07137_ _07139_ _07207_ _07208_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__or4_1
XANTENNA__12995__A2 _07455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15869__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ net1302 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_125_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11665_ _06324_ _06489_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__xnor2_1
X_14453_ net1276 vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17275__1334 vssd1 vssd1 vccd1 vccd1 _17275__1334/HI net1334 sky130_fd_sc_hd__conb_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10616_ _06146_ _06153_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__nand2_1
X_13404_ team_04_WB.MEM_SIZE_REG_REG\[19\] _07746_ _07829_ vssd1 vssd1 vccd1 vccd1
+ _07830_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12747__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_X net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17172_ clknet_leaf_92_wb_clk_i _02784_ _01401_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_14384_ net1457 vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_output190_A net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11596_ net532 _07046_ _07084_ net556 vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__a211o_1
XANTENNA__12009__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ net1086 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 _07761_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16123_ clknet_leaf_92_wb_clk_i _01792_ _00352_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ _06103_ net1583 net1020 vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14505__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13266_ net70 net2649 net977 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__mux2_1
X_16054_ clknet_leaf_18_wb_clk_i _01723_ _00283_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03529_
+ _06053_ _06056_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a31o_1
XANTENNA__08503__A _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10752__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ net229 net649 vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__and2_1
XANTENNA__13172__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15005_ net1154 vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__inv_2
X_13197_ _03635_ net271 net999 _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__a22o_1
XANTENNA__12025__A net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__A0 _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A1 _04166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ net253 net2385 net511 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
XANTENNA__11864__A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ net2190 net352 _07494_ net440 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16956_ clknet_leaf_125_wb_clk_i _02625_ _01185_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12132__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ clknet_leaf_11_wb_clk_i _01584_ _00134_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_139_Right_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16887_ clknet_leaf_173_wb_clk_i _02556_ _01116_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[860\]
+ sky130_fd_sc_hd__dfrtp_1
X_15838_ clknet_leaf_90_wb_clk_i _01515_ _00065_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11870__Y _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ net1289 vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XANTENNA__12435__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08310_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__mux2_1
XANTENNA__12986__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09290_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\]
+ net858 vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08241_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_14 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1082 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_25 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12738__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08172_ net752 _03782_ _03726_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_95_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11946__B1 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10943__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__11758__B net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput121 net121 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput132 net132 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xoutput143 net143 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_140_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput154 net154 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12371__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput165 net165 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput176 net176 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput187 net187 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XANTENNA__12910__A2 net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput198 net198 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XANTENNA_fanout486_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07956_ _03560_ _03561_ _03565_ _03566_ net787 net809 vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09214__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__B net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07887_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\] vssd1 vssd1
+ vccd1 vccd1 _03502_ sky130_fd_sc_hd__inv_2
XANTENNA__08878__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13871__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout653_A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10685__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[963\]
+ net890 vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout820_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12809__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08725__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08508_ _04115_ _04116_ _04117_ _04118_ net824 net742 vssd1 vssd1 vccd1 vccd1 _04119_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09488_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08439_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[568\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12729__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _04439_ net636 _04557_ net635 net545 net537 vssd1 vssd1 vccd1 vccd1 _06939_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ net283 _05983_ _05984_ _05980_ net1058 vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11949__A _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12544__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _06766_ _06869_ net538 vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13120_ _07552_ net380 net300 net1844 vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _05630_ _05922_ _05923_ net623 net279 vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13154__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ _07512_ net376 net308 net1673 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a22o_1
X_10263_ net620 _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__nor2_1
XANTENNA__12362__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09453__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net2538 net516 _07454_ net445 vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a22o_1
XANTENNA__12901__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _05798_ _05801_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\]
+ net1075 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__o2bb2a_1
X_16810_ clknet_leaf_160_wb_clk_i _02479_ _01039_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08469__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout370 net372 vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_2
Xfanout381 _07679_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_2
X_16741_ clknet_leaf_4_wb_clk_i _02410_ _00970_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[714\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout392 _07672_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_6
XANTENNA__11468__A2 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13953_ net1564 net1069 _03310_ net264 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a22o_1
XANTENNA__14995__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10676__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ _07606_ net346 net387 net2493 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__a22o_1
X_16672_ clknet_leaf_139_wb_clk_i _02341_ _00901_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _02921_ _03261_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15623_ net1139 vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12835_ _07533_ net326 net392 net1800 vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a22o_1
XANTENNA__12417__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output203_A net203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15554_ net1219 vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__inv_2
X_12766_ _07493_ net327 net396 net1720 vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14505_ net1263 vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__inv_2
X_11717_ _06900_ _06902_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__xnor2_1
X_15485_ net1155 vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__inv_2
X_12697_ net2221 net405 net334 _07284_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ net1430 _02834_ _01475_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_42_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__inv_2
X_14436_ net1292 vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__inv_2
Xinput12 DAT_I[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11928__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 DAT_I[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 gpio_in[9] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_1
Xinput45 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_1
X_17155_ clknet_leaf_82_wb_clk_i net1298 _01384_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14367_ net1441 vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__clkbuf_1
X_11579_ _05194_ net365 _07066_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__o211a_1
XANTENNA__10763__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput56 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput67 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_1
Xhold807 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[328\] vssd1 vssd1
+ vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xinput78 wbs_dat_i[18] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_1
X_16106_ clknet_leaf_163_wb_clk_i _01775_ _00335_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_13318_ net1084 team_04_WB.MEM_SIZE_REG_REG\[20\] vssd1 vssd1 vccd1 vccd1 _07744_
+ sky130_fd_sc_hd__nor2_1
Xinput89 wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_1
Xhold818 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\] vssd1 vssd1
+ vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
X_17086_ clknet_leaf_76_wb_clk_i net2310 _01315_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_14298_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\] _03463_
+ net818 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__o21ai_1
Xhold829 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\] vssd1 vssd1
+ vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09349__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13145__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ clknet_leaf_6_wb_clk_i _01706_ _00266_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249_ net88 team_04_WB.ADDR_START_VAL_REG\[27\] net976 vssd1 vssd1 vccd1 vccd1
+ _01657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11156__A1 _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08790_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[786\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__mux2_1
XANTENNA__08379__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13499__A1_N net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16939_ clknet_leaf_15_wb_clk_i _02608_ _01168_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10667__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__A _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_146_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10003__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _05018_ _05019_ _05020_ _05021_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05022_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ _04949_ _04950_ _04951_ _04952_ net836 net749 vssd1 vssd1 vccd1 vccd1 _04953_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_138_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12959__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11092__A0 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A2 _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09273_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[937\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08183__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08224_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[29\] team_04_WB.instance_to_wrap.CPU_DAT_O\[29\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13968__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08155_ _03762_ _03763_ _03764_ _03765_ net792 net802 vssd1 vssd1 vccd1 vccd1 _03766_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout401_A _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12364__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_151_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12592__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08143__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13136__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13984__A _04583_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__X _05137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15972__Q team_04_WB.ADDR_START_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\]
+ net968 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__mux2_1
X_17274__1333 vssd1 vssd1 vccd1 vccd1 _17274__1333/HI net1333 sky130_fd_sc_hd__conb_1
XANTENNA__13208__B _06145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] net973 _03549_ vssd1 vssd1 vccd1
+ vccd1 _03550_ sky130_fd_sc_hd__o21a_4
XANTENNA__12112__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_X net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10658__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15704__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _04920_ _06438_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_127_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09609_ team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] net974 vssd1 vssd1 vccd1 vccd1
+ _05220_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10881_ net634 _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12539__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10848__A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input101_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12620_ net699 _06198_ _07590_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__or3_4
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12551_ net2165 net222 net422 vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11502_ _06978_ _06979_ _06984_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15270_ net1104 vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__inv_2
X_12482_ net608 net221 net683 vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14221_ team_04_WB.instance_to_wrap.final_design.uart.receiving net34 vssd1 vssd1
+ vccd1 vccd1 _03418_ sky130_fd_sc_hd__nor2_1
X_11433_ _06802_ _06921_ net559 vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__mux2_1
XANTENNA__11386__A1 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12583__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] vssd1 vssd1
+ vccd1 vccd1 _03372_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11364_ _04273_ _04301_ net360 vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _05532_ vssd1
+ vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__nor2_1
X_13103_ _07535_ net373 net299 net1875 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a22o_1
XANTENNA__13127__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14083_ net1485 _06112_ net1032 vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__mux2_1
X_11295_ _06782_ _06783_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__and2_1
XFILLER_0_131_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ _07495_ net367 net306 net1659 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a22o_1
X_10246_ _05564_ _05566_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nand2_1
XANTENNA__11689__A2 _06248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1110 net1115 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
Xfanout1121 net1123 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
Xfanout1132 net1135 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_4
XANTENNA__10522__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ net643 _03836_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1143 net1144 vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 net1156 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__buf_4
Xfanout1176 net1181 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_2
Xfanout1187 net1194 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__clkbuf_4
X_14985_ net1132 vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__inv_2
Xfanout1198 net1202 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__buf_2
XFILLER_0_92_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16724_ clknet_leaf_3_wb_clk_i _02393_ _00953_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\]
+ sky130_fd_sc_hd__dfrtp_1
X_13936_ net1900 net1073 net1040 _03300_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10113__A2 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__X _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16655_ clknet_leaf_188_wb_clk_i _02324_ _00884_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13867_ _02897_ _03222_ _03223_ net1039 vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_9_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15606_ net1228 vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12818_ net232 net2288 net324 vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__mux2_1
X_16586_ clknet_leaf_160_wb_clk_i _02255_ _00815_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\]
+ sky130_fd_sc_hd__dfrtp_1
X_13798_ net998 _03185_ _03188_ _03183_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11074__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15537_ net1272 vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12749_ _07474_ net343 net402 net2101 vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10821__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15468_ net1121 vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__inv_2
X_17207_ net1413 _02817_ _01441_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_14419_ net1275 vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15399_ net1139 vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12574__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17138_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[3\]
+ _01367_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_163_1148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold604 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\] vssd1 vssd1
+ vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\] vssd1 vssd1
+ vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\] vssd1 vssd1
+ vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13118__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold637 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\] vssd1 vssd1
+ vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\] vssd1 vssd1
+ vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap356 _06600_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__buf_1
X_17069_ clknet_leaf_48_wb_clk_i _00016_ _01298_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_09960_ net591 _04387_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold659 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\] vssd1 vssd1
+ vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10780__X _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09493__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
X_09891_ _05499_ _05501_ _04303_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_0_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08842_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__mux2_1
X_08773_ net765 _04377_ _04383_ _04371_ vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11837__C1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11771__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11852__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout351_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout449_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_101_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09325_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1260_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout616_A _06192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09256_ net630 _04865_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__xor2_1
XANTENNA__08572__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15967__Q team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08207_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__mux2_1
XANTENNA__09105__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09187_ _04794_ _04795_ _04796_ _04797_ net824 net733 vssd1 vssd1 vccd1 vccd1 _04798_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_90_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_170_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_X net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__B2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08138_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13109__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _03676_ _03677_ _03678_ _03679_ net827 net735 vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12822__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _03499_ _04839_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2_1
XANTENNA__08023__D _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ net547 _05404_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ _05568_ _05640_ _05570_ _05567_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ net1238 vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11982_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _05342_ vssd1
+ vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__xor2_1
X_13721_ _07805_ _07811_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09432__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _06418_ _06420_ _06397_ _06400_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__a211o_1
XANTENNA__10578__A team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ clknet_leaf_151_wb_clk_i _02109_ _00669_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\]
+ sky130_fd_sc_hd__dfrtp_1
X_13652_ team_04_WB.ADDR_START_VAL_REG\[4\] _03042_ vssd1 vssd1 vccd1 vccd1 _03043_
+ sky130_fd_sc_hd__and2_1
X_10864_ net638 _06351_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__nor2_1
XANTENNA__13045__A1 _07506_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _07572_ net484 net413 net1815 vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16371_ clknet_leaf_182_wb_clk_i _02040_ _00600_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\]
+ sky130_fd_sc_hd__dfrtp_1
X_13583_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] net1044 _02973_
+ net1081 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ _06269_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15322_ net1146 vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__inv_2
XANTENNA__08472__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12534_ net2547 net260 net421 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08335__X _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15877__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15253_ net1207 vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__inv_2
XANTENNA__10517__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ net522 net602 _07466_ net429 net1966 vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a32o_1
XANTENNA__11359__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14204_ _03519_ _03407_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__nor2_1
XANTENNA__08224__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _06432_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__xor2_1
XANTENNA__12020__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15184_ net1160 vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__inv_2
X_12396_ net653 net607 net214 vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12017__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ net1090 net1088 net1089 net1087 vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11347_ _04087_ net363 vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14513__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14066_ net1446 _06078_ net1033 vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__mux2_1
X_11278_ net639 _04328_ net591 _04439_ net544 net535 vssd1 vssd1 vccd1 vccd1 _06767_
+ sky130_fd_sc_hd__mux4_2
XANTENNA__10760__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__xnor2_1
X_13017_ _07652_ net473 net312 net2030 vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a22o_1
XANTENNA__12033__A _07380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11531__A1 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net162 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_85_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12087__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14968_ net1222 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__inv_2
XANTENNA__08657__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16707_ clknet_leaf_125_wb_clk_i _02376_ _00936_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11591__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ _03118_ _03288_ _03110_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11834__A2 _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14899_ net1237 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10919__C net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16638_ clknet_leaf_129_wb_clk_i _02307_ _00867_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_162_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13799__A team_04_WB.ADDR_START_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16569_ clknet_leaf_152_wb_clk_i _02238_ _00798_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ _04717_ _04718_ _04719_ _04720_ net792 net815 vssd1 vssd1 vccd1 vccd1 _04721_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09488__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17273__1332 vssd1 vssd1 vccd1 vccd1 _17273__1332/HI net1332 sky130_fd_sc_hd__conb_1
XFILLER_0_142_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11112__A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold401 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\] vssd1 vssd1
+ vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold412 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[312\] vssd1 vssd1
+ vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\] vssd1 vssd1
+ vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 net128 vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10951__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold456 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\] vssd1 vssd1
+ vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\] vssd1 vssd1
+ vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\] vssd1 vssd1
+ vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09943_ net642 net660 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__nor2_1
Xhold489 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\] vssd1 vssd1
+ vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_61_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout903 net904 vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net926 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__clkbuf_4
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__buf_2
Xfanout936 net937 vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout399_A _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_161_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_161_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout947 net950 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_4
X_09874_ _05481_ _05482_ _05484_ _04979_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_146_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout958 net962 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_146_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout969 net970 vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__clkbuf_4
Xhold1101 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\] vssd1 vssd1
+ vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\] vssd1 vssd1
+ vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__mux2_1
Xhold1123 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\] vssd1 vssd1
+ vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\] vssd1 vssd1
+ vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[915\] vssd1 vssd1
+ vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\] vssd1 vssd1
+ vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\] vssd1 vssd1
+ vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__mux2_1
Xhold1178 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\] vssd1 vssd1
+ vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1189 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[352\] vssd1 vssd1
+ vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout733_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _04292_ _04297_ net720 vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__A1 _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1263_X net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09308_ net667 _04918_ _04894_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a21oi_2
X_10580_ _06125_ net1557 net1023 vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13996__X _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09239_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11022__A team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ _07320_ net672 vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout890_X net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__A1 _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ net558 _06689_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ net236 net647 vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__and2_1
XANTENNA__12552__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11132_ _06615_ _06620_ net576 vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold990 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\] vssd1 vssd1
+ vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
X_15940_ clknet_leaf_52_wb_clk_i _01617_ _00167_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__dfrtp_1
X_11063_ net592 net543 _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11513__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _05593_ _05624_ _05594_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12710__B1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ clknet_leaf_86_wb_clk_i _01548_ _00098_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_14822_ net1108 vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12069__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14753_ net1149 vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ net691 _07102_ _07425_ net614 vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__o211a_2
XANTENNA__08142__A0 _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13704_ team_04_WB.ADDR_START_VAL_REG\[7\] _02999_ _03002_ _03004_ vssd1 vssd1 vccd1
+ vccd1 _03095_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_80_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10916_ net565 _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_106_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14684_ net1126 vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11896_ net687 _07364_ _07365_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__a211o_1
XANTENNA__09890__B1 _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09317__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16423_ clknet_leaf_24_wb_clk_i _02092_ _00652_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\]
+ sky130_fd_sc_hd__dfrtp_1
X_13635_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] net1059 net1101
+ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ net596 _06335_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12777__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16354_ clknet_leaf_140_wb_clk_i _02023_ _00583_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13566_ team_04_WB.ADDR_START_VAL_REG\[15\] _02955_ vssd1 vssd1 vccd1 vccd1 _02957_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12241__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10778_ net583 net569 net466 _06202_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_4_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09101__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15305_ net1137 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12517_ _07514_ net490 net427 net1773 vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16285_ clknet_leaf_129_wb_clk_i _01954_ _00514_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _07733_ _07854_ _07857_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15236_ net1189 vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ net605 net218 net685 vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09608__Y _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ net1250 vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12379_ net243 net2550 net495 vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XANTENNA__11752__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_14118_ team_04_WB.MEM_SIZE_REG_REG\[17\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[17\]
+ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__a22o_1
XFILLER_0_120_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ net1151 vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14049_ net7 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1
+ vccd1 vccd1 _01537_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__B1 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09771__S net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_145_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4__f_wb_clk_i_A clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[436\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15074__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__mux2_1
XANTENNA__13257__A1 team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13306__B team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08541_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[54\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__mux2_1
XANTENNA__13009__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ net661 _04081_ _04082_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_106_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10011__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10946__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12768__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout314_A _07677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1056_A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[622\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13976__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold220 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\] vssd1 vssd1
+ vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13732__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12225__X _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 net150 vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_184_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold242 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\] vssd1 vssd1
+ vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold253 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\] vssd1 vssd1
+ vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold264 team_04_WB.instance_to_wrap.final_design.uart.working_data\[5\] vssd1 vssd1
+ vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[33\] vssd1 vssd1
+ vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout700 _05222_ vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__clkbuf_2
Xhold286 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\] vssd1 vssd1
+ vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\] vssd1 vssd1
+ vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13992__A _04811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09926_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _05536_ vssd1
+ vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout733 net736 vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__buf_4
Xfanout744 net750 vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
Xfanout755 _03626_ vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09681__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout766 net769 vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__buf_6
X_09857_ _04669_ _04726_ _05466_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout850_A net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout777 _03564_ vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__clkbuf_8
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 _03559_ vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__buf_4
XANTENNA__13056__X _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _04415_ _04416_ _04417_ _04418_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04419_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13248__A1 team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08297__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\]
+ net960 vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__mux2_1
X_08739_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[787\]
+ net870 vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
XANTENNA__12120__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15803__22 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__inv_2
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15712__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ _05451_ _06200_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__and3_2
XFILLER_0_138_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12471__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08029__C _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _04782_ _05279_ net822 vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__or3_1
XFILLER_0_166_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10482__B2 team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11681_ team_04_WB.MEM_SIZE_REG_REG\[23\] _06513_ vssd1 vssd1 vccd1 vccd1 _07170_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__12547__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_X net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ _07743_ _07845_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__nor2_1
X_10632_ _06162_ _06163_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__or3_1
XFILLER_0_165_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _07775_ _07776_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__nor2_1
XANTENNA__11431__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] net1095 net1051 vssd1 vssd1 vccd1
+ vccd1 _06114_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13971__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ net1916 net499 _07595_ net441 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070_ clknet_leaf_19_wb_clk_i _01739_ _00299_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10494_ _06046_ _06067_ _06068_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__o21ai_1
XANTENNA_input77_A wbs_dat_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] _07712_ _05525_
+ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13184__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15021_ net1152 vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ net2356 net505 _07559_ net452 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__a22o_1
X_12164_ net1989 net507 _07523_ net450 vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08061__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ _06222_ _06230_ net537 vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__mux2_1
X_16972_ clknet_leaf_112_wb_clk_i _02641_ _01201_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\]
+ sky130_fd_sc_hd__dfrtp_1
X_12095_ net2588 net355 _07502_ net458 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__a22o_1
XANTENNA__09591__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15923_ clknet_leaf_70_wb_clk_i _01600_ _00150_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11693__Y _07182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11046_ _06532_ _06534_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09786__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ clknet_leaf_95_wb_clk_i _01531_ _00081_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14805_ net1200 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08115__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ _07646_ net468 net310 net2267 vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a22o_1
XANTENNA__12998__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14736_ net1165 vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11948_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[5\] team_04_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ _07234_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08210__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14667_ net1167 vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__inv_2
X_11879_ _03613_ _05904_ _06184_ _04559_ net694 vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16406_ clknet_leaf_10_wb_clk_i _02075_ _00635_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\]
+ sky130_fd_sc_hd__dfrtp_1
X_13618_ _07691_ _03008_ net995 vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__a21o_1
XANTENNA__08418__A1 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12214__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14598_ net1185 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16337_ clknet_leaf_180_wb_clk_i _02006_ _00566_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _02937_ _02939_ net997 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10776__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16268_ clknet_leaf_111_wb_clk_i _01937_ _00497_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[241\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13175__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ net1233 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__inv_2
XANTENNA__15069__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16199_ clknet_leaf_24_wb_clk_i _01868_ _00428_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08277__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12205__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14124__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07972_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[735\]
+ net934 vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09711_ _05318_ _05319_ _05320_ _05321_ net797 net817 vssd1 vssd1 vccd1 vccd1 _05322_
+ sky130_fd_sc_hd__mux4_1
X_09642_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__mux2_1
XANTENNA__12221__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09573_ _05180_ _05181_ _05182_ _05183_ net833 net745 vssd1 vssd1 vccd1 vccd1 _05184_
+ sky130_fd_sc_hd__mux4_1
X_08524_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[951\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12453__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08845__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[88\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_1
XANTENNA__12367__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout431_A _07641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1173_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _06195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08386_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__mux2_1
XANTENNA__13402__A1 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09676__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13166__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ net1008 net1007 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[462\]
+ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_167_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12913__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15788__7 clknet_leaf_66_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__inv_2
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout530 net531 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14130__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _05518_ _05519_ _05470_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__mux2_1
Xfanout552 _05376_ vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
Xfanout563 net565 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_2
Xfanout585 net587 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__buf_2
X_12920_ _07622_ net344 net386 net1813 vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__a22o_1
Xfanout596 _04055_ vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__buf_2
XANTENNA__11673__C net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12692__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ _07549_ net341 net394 net1914 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_9__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__11970__A _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ net704 _05818_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__nor2_1
X_15570_ net1245 vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_3__f_wb_clk_i_X clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08755__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12782_ _07509_ net343 net398 net1651 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14521_ net1186 vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11733_ _07220_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12995__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ net1301 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14452_ net1278 vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _07151_ _07152_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_25_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10207__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ _07750_ _07825_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10615_ net58 _06152_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and2b_1
X_17171_ clknet_leaf_92_wb_clk_i _02783_ _01400_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13944__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14383_ net1443 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ _06568_ _06572_ net532 vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11955__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16122_ clknet_leaf_40_wb_clk_i _01791_ _00351_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07895__A team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09586__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13334_ net1086 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 _07760_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[18\]
+ _06102_ net1047 vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output183_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13157__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ clknet_leaf_33_wb_clk_i _01722_ _00282_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_13265_ net71 team_04_WB.ADDR_START_VAL_REG\[11\] net977 vssd1 vssd1 vccd1 vccd1
+ _01641_ sky130_fd_sc_hd__mux2_1
XANTENNA__10525__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_94_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10477_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] net1006 _06048_ _06052_
+ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11707__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ net1130 vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__inv_2
XANTENNA__12904__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__B2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ net1951 net509 _07549_ net451 vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a22o_1
X_13196_ net992 net991 vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12025__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12147_ net254 net2347 net512 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XANTENNA__14521__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14121__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__B _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ net248 net677 vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__and2_1
X_16955_ clknet_leaf_97_wb_clk_i _02624_ _01184_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[928\]
+ sky130_fd_sc_hd__dfrtp_1
X_11029_ team_04_WB.MEM_SIZE_REG_REG\[30\] team_04_WB.MEM_SIZE_REG_REG\[29\] _06517_
+ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__or3_1
X_15906_ clknet_leaf_36_wb_clk_i _01583_ _00133_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08431__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16886_ clknet_leaf_14_wb_clk_i _02555_ _01115_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\]
+ sky130_fd_sc_hd__dfrtp_1
X_15837_ clknet_leaf_91_wb_clk_i _01514_ _00064_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13571__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15768_ net1289 vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__inv_2
XANTENNA__12435__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14719_ net1241 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__inv_2
X_15794__13 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__inv_2
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15699_ net1268 vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[989\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_26 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_37 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[28\] team_04_WB.instance_to_wrap.CPU_DAT_O\[28\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__mux2_2
XFILLER_0_7_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17279__A net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10783__X _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09496__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13148__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput122 net122 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput133 net133 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput144 net144 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput155 net155 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput166 net166 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
Xoutput177 net177 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput188 net188 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput199 net199 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_162_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09084__X _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14112__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_07955_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout381_A _07679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08878__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07886_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\] vssd1
+ vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__inv_2
X_09625_ net724 _05229_ net714 vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10685__B2 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1290_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A _03589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09556_ _03724_ _04002_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__nand2_1
XANTENNA__13623__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08507_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[439\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08725__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ net774 _05091_ _05097_ net763 vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout813_A net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08438_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[632\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[600\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_156_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13926__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire216 _07264_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_2
X_08369_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[505\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[473\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11937__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire238 _07313_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__buf_2
X_10400_ net617 _05981_ net283 vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11380_ net636 _04557_ net546 vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__mux2_1
XANTENNA__11401__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _05708_ _05752_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10572__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10262_ _05763_ _05861_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or2_1
X_13050_ _07511_ net378 net308 net1627 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12001_ net217 net681 vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__and2_1
XANTENNA__08042__C net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ net281 _05800_ net1058 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08030__A2 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14103__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout360 _06254_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
Xfanout371 net372 vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_4
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16740_ clknet_leaf_169_wb_clk_i _02409_ _00969_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout382 net383 vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__clkbuf_4
Xfanout393 _07672_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_4
X_13952_ _03752_ net599 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__and2b_1
XANTENNA__13862__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ _07605_ net335 net385 net2185 vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22o_1
XANTENNA__10676__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16671_ clknet_leaf_157_wb_clk_i _02340_ _00900_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[644\]
+ sky130_fd_sc_hd__dfrtp_1
X_13883_ net2609 net1068 _03264_ _03265_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15622_ net1103 vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__inv_2
XANTENNA__15172__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ _07532_ net326 net392 net2136 vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12417__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15553_ net1129 vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12765_ _07492_ net329 net396 net1840 vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__a22o_1
XANTENNA__12968__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08057__Y _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13090__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14504_ net1259 vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__inv_2
X_11716_ _06782_ _06783_ _06918_ _07203_ _07204_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_84_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15484_ net1127 vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__inv_2
X_12696_ net2199 net405 net333 _07278_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17223_ net1429 _02833_ _01473_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14435_ net1292 vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _07040_ _07135_ _07077_ _07059_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_25_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11928__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 DAT_I[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ clknet_leaf_84_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[8\]
+ _01383_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput24 DAT_I[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 wb_rst_i vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_4
X_14366_ net1447 vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__clkbuf_1
Xinput46 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_1
XFILLER_0_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11578_ _05166_ _05192_ net361 vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__a21o_1
Xinput57 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_1
XFILLER_0_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput68 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_1
XFILLER_0_123_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16105_ clknet_leaf_121_wb_clk_i _01774_ _00334_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_13317_ team_04_WB.MEM_SIZE_REG_REG\[22\] _07741_ _07742_ vssd1 vssd1 vccd1 vccd1
+ _07743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold808 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\] vssd1 vssd1
+ vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput79 wbs_dat_i[19] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_1
X_17085_ clknet_leaf_76_wb_clk_i net1606 _01314_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10529_ _06091_ net1772 net1022 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold819 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\] vssd1 vssd1
+ vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_172_Right_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14297_ _03463_ _03464_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ clknet_leaf_20_wb_clk_i _01705_ _00265_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13248_ net89 team_04_WB.ADDR_START_VAL_REG\[28\] net976 vssd1 vssd1 vccd1 vccd1
+ _01658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11875__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _07615_ net380 net293 net1911 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a22o_1
XANTENNA__11594__B _07082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16938_ clknet_leaf_166_wb_clk_i _02607_ _01167_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10667__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_16869_ clknet_leaf_170_wb_clk_i _02538_ _01098_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\]
+ sky130_fd_sc_hd__dfrtp_1
X_09410_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[935\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08395__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09809__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09341_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_138_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_186_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_186_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11092__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09272_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[969\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_62_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_115_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _03816_ _03822_ _03833_ net767 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a22o_4
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout227_A _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08154_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[28\]
+ net950 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_151_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08085_ net646 _03694_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__xor2_4
XFILLER_0_113_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout596_A _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12344__B2 net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__B net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12380__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08643__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout763_A net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ net776 _04591_ net764 vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[17\] net1010
+ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__or2_1
XANTENNA__12647__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10658__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_X net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout649_X net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ net767 _05218_ _05207_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _04697_ _06295_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_973 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11607__A0 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09539_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[101\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[69\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__mux2_1
X_17289__1345 vssd1 vssd1 vccd1 vccd1 _17289__1345/HI net1345 sky130_fd_sc_hd__conb_1
XFILLER_0_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11025__A team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_159_Left_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12550_ net2507 net229 net422 vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11501_ _06699_ _06989_ _05139_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14021__A1 _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12481_ net2321 net430 _07653_ net524 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14336__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10864__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14220_ net1589 _06051_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11432_ _04328_ net591 _04439_ net636 net543 net536 vssd1 vssd1 vccd1 vccd1 _06921_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _03530_
+ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor3_1
XANTENNA__13780__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11363_ net567 _06602_ _06846_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13102_ _07534_ net373 net299 net1725 vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a22o_1
X_10314_ _05633_ _05906_ _05907_ net623 net279 vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14082_ net1496 _06110_ net1032 vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__mux2_1
X_11294_ net707 _06781_ _06762_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_168_Left_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13033_ _07494_ net371 net307 net1625 vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__a22o_1
X_10245_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] net1055 _05843_
+ _05846_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__a22o_1
XANTENNA__09200__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\] vssd1
+ vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12886__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1111 net1114 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__buf_4
X_10176_ net2647 net1058 _05782_ _05785_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a22o_1
Xfanout1122 net1123 vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
Xfanout1133 net1135 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__buf_2
Xfanout1144 net1157 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12303__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1155 net1156 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
Xfanout1166 net1187 vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__clkbuf_4
Xfanout1177 net1180 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
X_14984_ net1116 vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12638__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1188 net1194 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
Xfanout1199 net1201 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_4
X_13935_ _03091_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__xnor2_1
X_16723_ clknet_leaf_184_wb_clk_i _02392_ _00952_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13415__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload5_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16654_ clknet_leaf_30_wb_clk_i _02323_ _00883_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\]
+ sky130_fd_sc_hd__dfrtp_1
X_13866_ net1039 _03251_ _03252_ net1066 net1566 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__a32o_1
XANTENNA__08509__A net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10758__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ net1215 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__inv_2
XANTENNA__09104__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ net223 net2281 net324 vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16585_ clknet_leaf_123_wb_clk_i _02254_ _00814_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[558\]
+ sky130_fd_sc_hd__dfrtp_1
X_13797_ net1002 _03187_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15536_ net1173 vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__A1 net665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ _07473_ net347 net403 net2076 vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15467_ net1161 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
X_12679_ net234 net2551 net477 vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ net1412 _02816_ _01439_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14418_ net1289 vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15398_ net1103 vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__inv_2
X_17137_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[2\]
+ _01366_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14349_ net1191 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold605 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\] vssd1 vssd1
+ vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[576\] vssd1 vssd1
+ vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\] vssd1 vssd1
+ vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\] vssd1 vssd1
+ vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17068_ clknet_leaf_48_wb_clk_i _00015_ _01297_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold649 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\] vssd1 vssd1
+ vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_51_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16019_ clknet_leaf_75_wb_clk_i _01694_ _00248_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12326__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08910_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[528\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ _04359_ _05500_ _04329_ _04357_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08625__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12877__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08841_ net739 _04446_ net726 vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__a21o_1
XANTENNA__13309__B team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12213__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08772_ net778 _04382_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or2_1
XANTENNA__12629__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__B1 _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09014__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout344_A net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15540__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09324_ net781 _04934_ net764 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11604__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_153_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09255_ net630 _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout511_A net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12375__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1253_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout609_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08206_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09105__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09186_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_170_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_160_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08137_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08068_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[63\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[31\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15983__Q team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout880_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07992__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10328__B1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12868__A2 net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _05568_ _05640_ _05570_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11981_ net2359 net528 net457 _07439_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a22o_1
XANTENNA__10859__A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13720_ _06955_ net274 vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__nor2_1
X_10932_ _06418_ _06420_ _06400_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a21o_1
XANTENNA__10578__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13651_ net1000 _03038_ _03041_ _03037_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__o211a_1
X_10863_ net638 _06351_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08048__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11056__A1 _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12602_ _07571_ net493 net415 net2291 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16370_ clknet_leaf_10_wb_clk_i _02039_ _00599_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\]
+ sky130_fd_sc_hd__dfrtp_1
X_13582_ _07819_ _02972_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08763__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10794_ net587 _05192_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10264__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15321_ net1248 vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12533_ net2342 net246 net420 vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08472__A2 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15252_ net1225 vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__inv_2
X_12464_ net521 net605 _07465_ net429 net1894 vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a32o_1
XFILLER_0_136_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14203_ _03404_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[2\]
+ sky130_fd_sc_hd__and3_1
X_11415_ _06435_ _06903_ _06434_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a21oi_1
X_15183_ net1196 vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__inv_2
X_12395_ net1985 net434 _07626_ net523 vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14134_ net1091 net1088 vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nor2_1
XANTENNA_input62_X net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _06825_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__or2_1
XFILLER_0_162_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15893__Q net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12308__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14065_ net1456 _06076_ net1033 vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__mux2_1
X_11277_ _04385_ net545 _06229_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12859__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13016_ _07651_ net472 net312 net1873 vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a22o_1
X_10228_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] net1055 _05829_
+ _05831_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12033__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10159_ _05674_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and2_1
Xhold2 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[15\] vssd1 vssd1 vccd1
+ vccd1 net1439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ net1231 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__inv_2
X_16706_ clknet_leaf_147_wb_clk_i _02375_ _00935_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[679\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13918_ _03110_ _03118_ _03288_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__or3_1
XANTENNA__12492__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11591__C _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14898_ net1238 vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13849_ _03232_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16637_ clknet_leaf_132_wb_clk_i _02306_ _00866_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13036__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15360__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16568_ clknet_leaf_145_wb_clk_i _02237_ _00797_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15519_ net1273 vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__inv_2
X_16499_ clknet_leaf_182_wb_clk_i _02168_ _00728_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[172\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\]
+ net939 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09099__S0 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13744__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12923__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_60 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14704__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08846__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\] vssd1 vssd1
+ vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\] vssd1 vssd1
+ vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_174_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold424 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[548\] vssd1 vssd1
+ vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[594\] vssd1 vssd1
+ vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold446 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\] vssd1 vssd1
+ vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold457 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[720\] vssd1 vssd1
+ vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\] vssd1 vssd1
+ vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09942_ _03892_ _03894_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold479 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[828\] vssd1 vssd1
+ vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout904 _03657_ vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__buf_4
X_17288__1344 vssd1 vssd1 vccd1 vccd1 _17288__1344/HI net1344 sky130_fd_sc_hd__conb_1
Xfanout915 net926 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__buf_2
Xfanout926 _03555_ vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout937 net941 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_2
X_09873_ _05031_ _05086_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nand3_1
Xfanout948 net949 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_A _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_146_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\] vssd1 vssd1
+ vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
X_08824_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__mux2_1
Xhold1113 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\] vssd1 vssd1
+ vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10730__A0 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1001_A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\] vssd1 vssd1
+ vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08848__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1135 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\] vssd1 vssd1
+ vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\] vssd1 vssd1
+ vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08755_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[242\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[210\]
+ net936 vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
Xhold1157 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\] vssd1 vssd1
+ vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1168 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\] vssd1 vssd1
+ vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A _07252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09023__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1179 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\] vssd1 vssd1
+ vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout559_A _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ _04293_ _04294_ _04295_ _04296_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04297_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13027__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout726_A _03668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_172_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09100__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ _04900_ _04906_ _04917_ net716 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a22o_2
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12118__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09169_ _03591_ net759 _03656_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11200_ net644 _03891_ net642 net640 net544 net535 vssd1 vssd1 vccd1 vccd1 _06689_
+ sky130_fd_sc_hd__mux4_1
X_12180_ net2064 net507 _07531_ net443 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _06619_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[972\] vssd1 vssd1
+ vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\] vssd1 vssd1
+ vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net638 net549 vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__and2_1
XANTENNA__09262__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _04947_ _04948_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__o21ba_1
XANTENNA__11973__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15870_ clknet_leaf_95_wb_clk_i _01547_ _00097_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__08758__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A DAT_I[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1111 vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14752_ net1213 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__inv_2
XANTENNA__11277__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _07398_ _07424_ _07423_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08142__A1 _03752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ _03018_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__or2_1
X_10915_ net548 net542 net659 vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a21oi_1
X_14683_ net1145 vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11895_ net760 _05920_ _06184_ _04728_ net695 vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__a221o_1
XANTENNA__13018__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13634_ net1059 net1101 vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and2_1
X_16422_ clknet_leaf_17_wb_clk_i _02091_ _00651_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[395\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09317__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10846_ _04083_ _06304_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16353_ clknet_leaf_133_wb_clk_i _02022_ _00582_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13565_ team_04_WB.ADDR_START_VAL_REG\[15\] _02955_ vssd1 vssd1 vccd1 vccd1 _02956_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10528__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ net530 _06265_ net557 vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_165_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15304_ net1118 vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12516_ _07513_ net489 net426 net2096 vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a22o_1
X_16284_ clknet_leaf_116_wb_clk_i _01953_ _00513_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[257\]
+ sky130_fd_sc_hd__dfrtp_1
X_13496_ _07197_ net273 _07697_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12529__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15235_ net1170 vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12447_ net2430 net430 _07644_ net523 vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XANTENNA__14524__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15166_ net1215 vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_2
X_12378_ net255 net2324 net497 vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14117_ team_04_WB.MEM_SIZE_REG_REG\[16\] net988 net981 team_04_WB.ADDR_START_VAL_REG\[16\]
+ net1005 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__o221a_1
XFILLER_0_10_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11329_ net753 _06729_ _06731_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15097_ net1248 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ net8 net1061 net1037 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1
+ vccd1 vccd1 _01538_ sky130_fd_sc_hd__o22a_1
XFILLER_0_157_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12331__X _07610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15999_ clknet_leaf_51_wb_clk_i _01675_ _00228_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_141_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08540_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[86\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_141_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ net751 net717 _03726_ net662 vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12768__A1 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13322__B team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_114_Left_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09023_ _04630_ _04631_ _04632_ _04633_ net836 net739 vssd1 vssd1 vccd1 vccd1 _04634_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_A _07680_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold210 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\] vssd1 vssd1
+ vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\] vssd1 vssd1
+ vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold232 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\] vssd1 vssd1
+ vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09696__A1_N net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\] vssd1 vssd1
+ vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold254 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\] vssd1 vssd1
+ vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _02723_ vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\] vssd1 vssd1
+ vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1216_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold287 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\] vssd1 vssd1
+ vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout701 _05221_ vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_2
X_09925_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\]
+ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__and3_1
Xhold298 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[310\] vssd1 vssd1
+ vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout712 _03675_ vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout723 _03668_ vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
XANTENNA__13992__B net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13496__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout734 net736 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_123_Left_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout745 net747 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
XANTENNA_fanout676_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_X net297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_2
XANTENNA__07990__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _05466_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__inv_2
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_8
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net782 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__buf_4
XANTENNA__08578__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout789 net790 vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09263__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[433\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_8__f_wb_clk_i clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_09787_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout843_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _04276_ _04277_ _04278_ _04279_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04280_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09872__A1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B2 _05166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10700_ net1057 _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__or2_2
XFILLER_0_95_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11680_ _07166_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08890__A1_N net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__A1 _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _06164_ _06165_ _06166_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__or4_1
XANTENNA__09085__C1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ _07770_ _07774_ _07773_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10562_ _06113_ net1789 net1020 vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13971__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13708__B1 _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ net219 net670 vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__and2_1
X_13281_ _05613_ _07711_ net617 _07440_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__a2bb2o_1
X_10493_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] net1006 _06066_ vssd1
+ vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14344__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13184__A1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15020_ net1119 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12232_ net215 net674 vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__and2_1
X_12163_ net212 net649 vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _06227_ _06602_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__nor2_1
XANTENNA__09725__X _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16971_ clknet_leaf_15_wb_clk_i _02640_ _01200_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[944\]
+ sky130_fd_sc_hd__dfrtp_1
X_12094_ net256 net679 vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15922_ clknet_leaf_72_wb_clk_i _01599_ _00149_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__dfrtp_1
X_11045_ net645 net557 vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__nor2_1
XANTENNA__12695__B1 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__A1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15853_ clknet_leaf_86_wb_clk_i _01530_ _00080_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12311__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ net1208 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12996_ net601 _07456_ net468 net310 net1652 vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11947_ net905 _03630_ _05972_ _05975_ net756 vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__o32a_1
X_14735_ net1140 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08210__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14519__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14666_ net1124 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11878_ net705 _05899_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17287__1343 vssd1 vssd1 vccd1 vccd1 _17287__1343/HI net1343 sky130_fd_sc_hd__conb_1
XFILLER_0_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13617_ _03500_ _05968_ net1101 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__mux2_1
X_16405_ clknet_leaf_34_wb_clk_i _02074_ _00634_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__inv_2
X_14597_ net1184 vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__inv_2
XANTENNA__12039__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13548_ net992 _02936_ _02938_ net989 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16336_ clknet_leaf_1_wb_clk_i _02005_ _00565_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08951__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11878__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16267_ clknet_leaf_16_wb_clk_i _01936_ _00496_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13479_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] _05800_ net1100
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10782__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13175__A1 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15218_ net1246 vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09348__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16198_ clknet_leaf_18_wb_clk_i _01867_ _00427_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08252__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08277__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15149_ net1199 vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__inv_2
XANTENNA__14124__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09782__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire644_A _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07971_ _03578_ _03579_ _03580_ _03581_ net787 net810 vssd1 vssd1 vccd1 vccd1 _03582_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_71_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09710_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09641_ net579 net570 vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12221__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09572_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[901\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08523_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[983\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11110__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08454_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[184\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09530__B net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09022__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13938__B1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08385_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\]
+ net910 vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A _07656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1166_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12610__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13479__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12383__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10692__A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09006_ _04614_ _04616_ net739 vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o21a_1
XANTENNA__08162__A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout793_A net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_131_Left_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09692__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout581_X net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _06197_ vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__clkbuf_4
Xfanout531 net534 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout679_X net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout542 _05434_ vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_2
X_09908_ _05495_ _05511_ _05516_ _05440_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a31oi_2
XANTENNA__12677__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_2
Xfanout564 net565 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout575 _05250_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_2
Xfanout586 net587 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_2
X_09839_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__inv_2
XANTENNA__08101__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _07548_ net342 net394 net1991 vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11801_ net2271 net527 net446 _07284_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a22o_1
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12781_ _07508_ net347 net399 net1833 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_Left_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ net1186 vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__inv_2
X_11732_ _06973_ _06974_ _06992_ _06994_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__o22a_1
XFILLER_0_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14451_ net1272 vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__inv_2
X_11663_ team_04_WB.MEM_SIZE_REG_REG\[14\] _06507_ vssd1 vssd1 vccd1 vccd1 _07152_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_153_Right_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ team_04_WB.MEM_SIZE_REG_REG\[18\] _07747_ _07827_ vssd1 vssd1 vccd1 vccd1
+ _07828_ sky130_fd_sc_hd__a21bo_1
X_10614_ _06149_ _06150_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__nor3_1
XFILLER_0_153_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17170_ clknet_leaf_91_wb_clk_i _02782_ _01399_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12601__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ net1501 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__clkbuf_1
X_11594_ _07081_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16121_ clknet_leaf_177_wb_clk_i _01790_ _00350_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13333_ _07757_ _07758_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net1095 net1051 vssd1 vssd1 vccd1
+ vccd1 _06102_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16052_ clknet_leaf_6_wb_clk_i _01721_ _00281_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_13264_ net72 team_04_WB.ADDR_START_VAL_REG\[12\] net977 vssd1 vssd1 vccd1 vccd1
+ _01642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10476_ _06028_ _06037_ _06043_ _06036_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or4b_1
XFILLER_0_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15003_ net1145 vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__inv_2
X_12215_ net231 net649 vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__and2_2
X_13195_ net1031 net1025 vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nand2_1
XANTENNA__10915__B1 net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09781__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ net243 net2404 net511 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09208__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14535__2 clknet_leaf_105_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__inv_2
XFILLER_0_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10541__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12668__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16954_ clknet_leaf_44_wb_clk_i _02623_ _01183_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\]
+ sky130_fd_sc_hd__dfrtp_1
X_12077_ net2253 net352 _07493_ net438 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XANTENNA__08336__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09107__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ team_04_WB.MEM_SIZE_REG_REG\[28\] _06516_ vssd1 vssd1 vccd1 vccd1 _06517_
+ sky130_fd_sc_hd__or2_2
X_15905_ clknet_leaf_124_wb_clk_i _01582_ _00132_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12041__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16885_ clknet_leaf_34_wb_clk_i _02554_ _01114_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08431__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15836_ clknet_leaf_93_wb_clk_i _01513_ _00063_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15767_ net1283 vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
XANTENNA__13093__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ net602 _07391_ net469 net314 net1932 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13632__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14718_ net1218 vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__inv_2
XANTENNA__12840__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15698_ net1268 vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14649_ net1241 vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__inv_2
XANTENNA_16 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_27 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09777__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ net767 _03773_ _03779_ _03761_ _03767_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__a32o_2
XTAP_TAPCELL_ROW_136_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11946__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16319_ clknet_leaf_155_wb_clk_i _01988_ _00548_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17299_ net1355 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_15_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput123 net123 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput134 net134 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12931__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput145 net145 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
Xoutput156 net156 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput167 net167 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
Xoutput178 net178 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__clkbuf_4
Xoutput189 net189 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08710__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12659__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[511\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12123__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] vssd1 vssd1 vccd1
+ vccd1 _03500_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ net730 _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__nor2_1
XANTENNA__10685__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09555_ net767 _05165_ _05154_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13084__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12378__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1283_A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _04218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__X _06624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[503\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11634__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ net780 _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or2_1
X_08437_ _04044_ _04045_ _04046_ _04047_ net785 net806 vssd1 vssd1 vccd1 vccd1 _04048_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13998__A _04972_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1071_X net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15790__9 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout806_A net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09687__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[281\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11937__A2 _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08299_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[827\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17271__1331 vssd1 vssd1 vccd1 vccd1 _17271__1331/HI net1331 sky130_fd_sc_hd__conb_1
X_10330_ _05587_ _05629_ net618 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_971 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09438__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ _05688_ _05762_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12898__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14622__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ net2362 net515 _07453_ net441 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a22o_1
XANTENNA__08042__D net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _05542_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17286__1342 vssd1 vssd1 vccd1 vccd1 _17286__1342/HI net1342 sky130_fd_sc_hd__conb_1
XANTENNA__10361__S net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_4
Xfanout361 _06254_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_2
Xfanout372 _07679_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_4
X_13951_ _03693_ net263 net598 _03306_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__a31o_1
Xfanout383 _07679_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_4
Xfanout394 _07672_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_8
X_12902_ _07604_ net339 net385 net1826 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__a22o_1
X_13882_ _02910_ _03263_ net1039 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__o21a_1
XANTENNA__10676__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16670_ clknet_leaf_142_wb_clk_i _02339_ _00899_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\]
+ sky130_fd_sc_hd__dfrtp_1
X_12833_ _07531_ net329 net392 net1842 vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__a22o_1
X_15621_ net1108 vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__inv_2
XANTENNA__13075__A0 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08177__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09170__B net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11625__A1 _06776_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12764_ _07491_ net327 net396 net1765 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a22o_1
X_15552_ net1212 vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14503_ net1285 vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__inv_2
X_11715_ _06816_ _06817_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15483_ net1136 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
X_12695_ net2239 net404 net330 _07272_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input92_X net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17222_ net1428 _02832_ _01471_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09597__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11646_ _07117_ _07131_ _07132_ _07134_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or4_1
X_14434_ net1291 vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput14 DAT_I[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
X_17153_ clknet_leaf_84_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[7\]
+ _01382_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput25 DAT_I[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
X_14365_ net1479 vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__clkbuf_1
Xinput36 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12050__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _05166_ _05192_ net359 vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__or3_1
XANTENNA__12317__A _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
Xinput58 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
X_13316_ _07738_ _07740_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__a21oi_1
X_16104_ clknet_leaf_113_wb_clk_i _01773_ _00333_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_161_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput69 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
X_17084_ clknet_leaf_43_wb_clk_i _00040_ _01313_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.receiving
+ sky130_fd_sc_hd__dfrtp_2
X_10528_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[24\]
+ _06090_ net1049 vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__mux2_1
X_14296_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] _03462_
+ net818 vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold809 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\] vssd1 vssd1
+ vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13247_ net90 team_04_WB.ADDR_START_VAL_REG\[29\] net976 vssd1 vssd1 vccd1 vccd1
+ _01659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_0_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16035_ clknet_leaf_117_wb_clk_i _01704_ _00264_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10459_ _06030_ _06034_ _06035_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13178_ _07614_ net372 net291 net1919 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a22o_1
XANTENNA__08530__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ net214 net2451 net513 vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XANTENNA__12105__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A0 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16937_ clknet_leaf_99_wb_clk_i _02606_ _01166_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08404__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10667__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16868_ clknet_leaf_173_wb_clk_i _02537_ _01097_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\]
+ sky130_fd_sc_hd__dfrtp_1
X_15819_ clknet_leaf_85_wb_clk_i _01496_ _00046_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ clknet_leaf_159_wb_clk_i _02468_ _01028_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09340_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[232\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__mux2_1
XANTENNA__12813__A0 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09271_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[777\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_726 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12926__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _03827_ _03832_ net774 vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11919__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13330__B team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[124\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\]
+ net946 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_155_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_155_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_151_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12592__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _03694_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__inv_2
XFILLER_0_113_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12661__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__A _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07982__C net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08643__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ net781 _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__nor2_1
X_07937_ _03540_ net1024 vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10658__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08720__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13057__A0 _07246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09607_ _05212_ _05217_ net775 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout923_A net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_805 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12804__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[133\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11607__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09469_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14617__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ net577 _06987_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12480_ net608 net229 net682 vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__and3_1
XANTENNA__09210__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11431_ _06454_ _06919_ net464 vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__B2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10043__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] vssd1 vssd1
+ vccd1 vccd1 _03370_ sky130_fd_sc_hd__o21a_1
XANTENNA__13780__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12583__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ net587 _06849_ _06850_ _06272_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11791__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ _07533_ net368 net298 net1666 vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ _05703_ _05754_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14081_ net1469 _06108_ net1032 vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ net707 _06781_ _06762_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__or3b_1
XFILLER_0_104_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14352__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ _07493_ net369 net306 net1795 vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__a22o_1
XANTENNA_input52_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ net277 _05845_ net1074 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__o21a_1
XANTENNA__09446__A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1102 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1112 net1114 vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_125_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ net281 _05784_ net1056 vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__a21oi_1
Xfanout1123 net1158 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_2
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__buf_4
Xfanout1145 net1147 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_4
Xfanout1156 net1157 vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_2
XFILLER_0_156_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1167 net1169 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__buf_4
X_14983_ net1139 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__inv_2
XANTENNA__12099__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1178 net1180 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
Xfanout1189 net1194 vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08398__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16722_ clknet_leaf_18_wb_clk_i _02391_ _00951_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\]
+ sky130_fd_sc_hd__dfrtp_1
X_13934_ _03043_ _03087_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__nor2_1
XANTENNA__11846__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ clknet_leaf_28_wb_clk_i _02322_ _00882_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[626\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13048__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13865_ _02895_ _03250_ _02886_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15604_ net1235 vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__inv_2
X_12816_ net233 net2409 net324 vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16584_ clknet_leaf_160_wb_clk_i _02253_ _00813_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13796_ net992 _03184_ _03186_ net990 vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ net1195 vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__inv_2
XANTENNA__11074__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12747_ _07472_ net330 net400 net1984 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__a22o_1
XANTENNA__14527__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12271__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10282__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10821__A2 _06308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ net261 net2528 net477 vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__mux2_1
X_15466_ net1107 vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09120__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17205_ net1411 _02815_ _01437_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_11629_ team_04_WB.MEM_SIZE_REG_REG\[3\] team_04_WB.MEM_SIZE_REG_REG\[2\] team_04_WB.MEM_SIZE_REG_REG\[4\]
+ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__a21oi_1
X_14417_ net1290 vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15397_ net1109 vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__inv_2
XANTENNA__12047__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17136_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[1\]
+ _01365_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12574__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ net1191 vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_164_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold606 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\] vssd1 vssd1
+ vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11782__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold617 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[313\] vssd1 vssd1
+ vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\] vssd1 vssd1
+ vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
X_17067_ clknet_leaf_48_wb_clk_i _00014_ _01296_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_14279_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[21\] _03452_
+ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__and2_1
Xhold639 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[456\] vssd1 vssd1
+ vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10790__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12326__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ clknet_leaf_83_wb_clk_i _00006_ _00247_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08625__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08840_ _04448_ _04450_ net748 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08771_ _04378_ _04379_ _04380_ _04381_ net789 net810 vssd1 vssd1 vccd1 vccd1 _04382_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13606__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15093__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11837__A1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270__1330 vssd1 vssd1 vccd1 vccd1 _17270__1330/HI net1330 sky130_fd_sc_hd__conb_1
XFILLER_0_149_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13039__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09323_ _04930_ _04931_ _04932_ _04933_ net796 net803 vssd1 vssd1 vccd1 vccd1 _04934_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12656__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout337_A _07667_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10273__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ net666 _04864_ _04840_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_146_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17285__1341 vssd1 vssd1 vccd1 vccd1 _17285__1341/HI net1341 sky130_fd_sc_hd__conb_1
XFILLER_0_69_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08205_ net774 _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__or2_1
XANTENNA__13211__A0 net92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12014__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout504_A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1246_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[830\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15268__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[95\]
+ net866 vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12391__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10328__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15__f_wb_clk_i_X clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__B net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout661_X net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11980_ net655 _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09205__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _06400_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10578__C net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13650_ net1000 _07693_ _03035_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nand4_1
X_10862_ _04300_ _06300_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _07570_ net486 net413 net1872 vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a22o_1
XANTENNA__08048__C net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13581_ _07767_ _07815_ _07766_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12253__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _04300_ net657 vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__nand2_1
XANTENNA__14347__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15320_ net1204 vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__inv_2
X_12532_ net2206 net236 net420 vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15251_ net1233 vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ _06197_ net610 _07464_ net431 net1760 vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__a32o_1
XFILLER_0_152_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14202_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1090
+ net1089 vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a21o_1
X_11414_ _06383_ _06427_ _06440_ _06446_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__a31o_1
XANTENNA__12556__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15182_ net1204 vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__inv_2
X_12394_ net653 net607 net212 vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__and3_1
XANTENNA__08632__X _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[9\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[8\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__or4_1
XFILLER_0_22_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ _06272_ _06833_ _06830_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12308__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14064_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\] net1077
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] vssd1 vssd1
+ vccd1 vccd1 _03354_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09176__A _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ net595 net593 net592 net638 net545 net535 vssd1 vssd1 vccd1 vccd1 _06765_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10319__B2 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ _07650_ net472 net312 net2049 vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_18_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10227_ net277 _05830_ net1074 vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13269__A0 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11531__A3 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _05675_ _05768_ _05676_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_33_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 net147 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11819__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ _04612_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] vssd1
+ vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__and2b_1
X_14966_ net1228 vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10769__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16705_ clknet_leaf_133_wb_clk_i _02374_ _00934_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\]
+ sky130_fd_sc_hd__dfrtp_1
X_13917_ _03144_ _03287_ _03121_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14897_ net1265 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16636_ clknet_leaf_126_wb_clk_i _02305_ _00865_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13848_ net998 _03238_ _03236_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08954__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16567_ clknet_leaf_175_wb_clk_i _02236_ _00796_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\]
+ sky130_fd_sc_hd__dfrtp_1
X_13779_ _03159_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_100_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11380__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15518_ net1216 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16498_ clknet_leaf_9_wb_clk_i _02167_ _00727_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15449_ net1251 vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09099__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08846__S1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\] vssd1 vssd1
+ vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17119_ clknet_leaf_67_wb_clk_i _02754_ _01348_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold414 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\] vssd1 vssd1
+ vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold425 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\] vssd1 vssd1
+ vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08620__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold436 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\] vssd1 vssd1
+ vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[383\] vssd1 vssd1
+ vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold458 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[120\] vssd1 vssd1
+ vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09941_ _03892_ _03894_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold469 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\] vssd1 vssd1
+ vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout905 _03607_ vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout916 net917 vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout927 net929 vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ net588 net583 _05194_ _05193_ _05166_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__a32o_1
Xfanout938 net939 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14720__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\] vssd1 vssd1
+ vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
X_08823_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\] vssd1 vssd1
+ vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09281__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10730__A1 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1125 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\] vssd1 vssd1
+ vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1136 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[280\] vssd1 vssd1
+ vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ net773 _04364_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or2_1
Xhold1147 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\] vssd1 vssd1
+ vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12240__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1158 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\] vssd1 vssd1
+ vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\] vssd1 vssd1
+ vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09023__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09025__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__mux2_1
XANTENNA__12483__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_A net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1196_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12386__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout621_A net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_170_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_170_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout719_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _04911_ _04916_ net721 vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__mux2_1
XANTENNA__09100__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12786__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09237_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09695__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09168_ net766 _04778_ _04767_ _04761_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__o2bb2a_2
XTAP_TAPCELL_ROW_118_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout990_A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\]
+ net851 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09099_ _04706_ _04707_ _04708_ _04709_ net798 net802 vssd1 vssd1 vccd1 vccd1 _04710_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _06616_ _06618_ net563 vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__mux2_1
XANTENNA__08104__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold970 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\] vssd1 vssd1
+ vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\] vssd1 vssd1
+ vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold992 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\] vssd1 vssd1
+ vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _06548_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__and2b_1
XANTENNA__09262__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ _05595_ _05621_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__o21a_1
XANTENNA__12710__A2 net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A3 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10721__A1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ net1169 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input15_A DAT_I[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751_ net1241 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__inv_2
XANTENNA__11277__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[3\] team_04_WB.instance_to_wrap.CPU_DAT_O\[3\]
+ net266 vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13702_ _03045_ _03086_ _03092_ _03090_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__o31a_1
XFILLER_0_6_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10914_ net579 _06402_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__nor2_1
X_11894_ net705 _05917_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__nor2_1
X_14682_ net1146 vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16421_ clknet_leaf_20_wb_clk_i _02090_ _00650_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13633_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] net1045 _03020_
+ net1098 vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__a2bb2o_1
X_10845_ net641 _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08525__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16352_ clknet_leaf_135_wb_clk_i _02021_ _00581_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12777__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13564_ net710 _02949_ _02951_ net998 _02954_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10776_ net645 net545 _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12309__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ net1142 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12515_ _07512_ net488 net426 net1832 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a22o_1
X_13495_ _02884_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__nor2_1
X_16283_ clknet_leaf_103_wb_clk_i _01952_ _00512_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[256\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13726__A1 _07696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13726__B2 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ net609 net219 net682 vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__and3_1
X_15234_ net1218 vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08362__X _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08803__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15165_ net1147 vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
X_12377_ net257 net2333 net498 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12325__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14116_ team_04_WB.MEM_SIZE_REG_REG\[15\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[15\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__o221a_1
X_11328_ team_04_WB.MEM_SIZE_REG_REG\[20\] _06511_ vssd1 vssd1 vccd1 vccd1 _06817_
+ sky130_fd_sc_hd__xor2_2
X_15096_ net1206 vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14047_ net9 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1
+ vccd1 vccd1 _01539_ sky130_fd_sc_hd__o22a_1
X_11259_ net585 _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nand2_1
XANTENNA__08949__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12701__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17284__1340 vssd1 vssd1 vccd1 vccd1 _17284__1340/HI net1340 sky130_fd_sc_hd__conb_1
XANTENNA__12060__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15998_ clknet_leaf_59_wb_clk_i _01674_ _00227_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_167_Right_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14949_ net1109 vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__inv_2
XANTENNA__12465__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08470_ _04063_ _04069_ _04080_ net716 vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__a22o_4
XANTENNA__09640__Y _05251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13009__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ clknet_leaf_30_wb_clk_i _02288_ _00848_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12768__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13965__A1 _04081_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11976__B1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12219__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12934__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09022_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[16\]
+ vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[0\] vssd1
+ vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold222 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\] vssd1 vssd1
+ vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold233 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\] vssd1 vssd1
+ vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10400__B1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[249\] vssd1 vssd1
+ vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold255 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[318\] vssd1 vssd1
+ vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold266 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\] vssd1 vssd1
+ vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold277 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\] vssd1 vssd1
+ vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[115\] vssd1 vssd1
+ vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05534_ vssd1
+ vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and2_1
Xfanout702 net703 vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__buf_4
Xhold299 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\] vssd1 vssd1
+ vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout713 _03675_ vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_4
XANTENNA__13992__C _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12153__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout735 net736 vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1209_A net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_165_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout746 net747 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_2
Xfanout757 _03614_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07990__C net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A DAT_I[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _04725_ _05444_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__and2_2
Xfanout768 net769 vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
Xfanout779 net782 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout669_A _07589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\]
+ net966 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__mux2_1
X_09786_ _05393_ _05394_ _05395_ _05396_ net794 net814 vssd1 vssd1 vccd1 vccd1 _05397_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08737_ _04344_ _04345_ _04346_ _04347_ net827 net735 vssd1 vssd1 vccd1 vccd1 _04348_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout457_X net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_A net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__A team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08668_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XANTENNA__10696__Y _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09872__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XANTENNA__12208__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10630_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[2\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\]
+ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__or4_1
XFILLER_0_154_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12759__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11967__B1 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[13\]
+ _06112_ net1047 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12300_ net2287 net501 _07594_ net450 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a22o_1
XANTENNA__13708__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ _05336_ _05341_ net617 vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__a21o_1
X_10492_ _06028_ _06045_ _06052_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12231_ net2531 net503 _07558_ net450 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13184__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ net2565 net508 _07522_ net448 vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11113_ net356 _06601_ net557 vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_9_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15456__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ net2242 net354 _07501_ net451 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a22o_1
X_16970_ clknet_leaf_162_wb_clk_i _02639_ _01199_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14360__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08769__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12144__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15921_ clknet_leaf_71_wb_clk_i _01598_ _00148_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09454__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ net645 net571 vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08363__A2 _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ clknet_leaf_86_wb_clk_i _01529_ _00079_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14803_ net1231 vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15783_ net1287 vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__inv_2
XANTENNA__12447__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10112__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12995_ net603 _07455_ net470 net311 net2260 vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14734_ net1198 vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__inv_2
XANTENNA__12998__A2 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946_ net2223 net528 net454 _07409_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14665_ net1132 vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__inv_2
X_11877_ net2335 net527 net446 _07350_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__a22o_1
X_16404_ clknet_leaf_2_wb_clk_i _02073_ _00633_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\]
+ sky130_fd_sc_hd__dfrtp_1
X_13616_ net993 _03006_ net999 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ net643 _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14596_ net1176 vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12039__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16335_ clknet_leaf_187_wb_clk_i _02004_ _00564_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13547_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] _05858_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__mux2_1
X_10759_ _05447_ net467 _05469_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__and3_4
XFILLER_0_70_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16266_ clknet_leaf_164_wb_clk_i _01935_ _00495_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13478_ net1002 _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10782__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13175__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15217_ net1271 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__inv_2
X_12429_ net2117 net434 _07635_ net524 vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16197_ clknet_leaf_5_wb_clk_i _01866_ _00426_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12383__A0 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15148_ net1128 vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13585__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11894__A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[927\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__mux2_1
XANTENNA__08679__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15079_ net1139 vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09364__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08985__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09640_ net664 _05248_ _05249_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__a21oi_2
Xclkbuf_leaf_109_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_160_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09571_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__mux2_1
XANTENNA__12929__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08522_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__mux2_1
XANTENNA__08737__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09303__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[248\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\]
+ net849 vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08384_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\]
+ net909 vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12664__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09005_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[302\] net899 net836
+ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__o211a_1
XANTENNA__13166__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12374__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09465__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12913__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout786_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14115__B2 team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout510 _07521_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__buf_4
Xfanout521 net522 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__clkbuf_4
X_09907_ _03696_ _05495_ _05511_ _05516_ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__a41oi_4
Xfanout532 net534 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__buf_2
Xfanout543 net544 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
XANTENNA_fanout953_A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 net556 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
Xfanout565 _05309_ vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
XANTENNA__10688__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
X_09838_ _05442_ _05446_ _05448_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__and3_1
Xfanout587 _05139_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
Xfanout598 net599 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12429__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _05336_ net551 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11800_ net652 net227 vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__and2_1
X_12780_ _07507_ net330 net396 net1751 vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a22o_1
XANTENNA__09213__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11101__B2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _06992_ _06994_ _06975_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10359__S net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14450_ net1276 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__inv_2
X_11662_ net707 _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _07746_ _07826_ _07747_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__o21bai_1
X_10613_ net60 net59 net56 net57 vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14381_ net1451 vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__clkbuf_1
X_11593_ _06743_ _06886_ _06948_ _06751_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14355__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16120_ clknet_leaf_153_wb_clk_i _01789_ _00349_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_13332_ team_04_WB.MEM_SIZE_REG_REG\[15\] _07756_ vssd1 vssd1 vccd1 vccd1 _07758_
+ sky130_fd_sc_hd__and2_1
XANTENNA_input82_A wbs_dat_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ _06101_ net1547 net1020 vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16051_ clknet_leaf_188_wb_clk_i _01720_ _00280_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13157__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ _06037_ _06043_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__or2_1
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13263_ net73 team_04_WB.ADDR_START_VAL_REG\[13\] net976 vssd1 vssd1 vccd1 vccd1
+ _01643_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_121_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12365__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15002_ net1152 vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__inv_2
XANTENNA__08033__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12214_ net2086 net509 _07548_ net453 vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a22o_1
XANTENNA__12904__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13194_ net1029 net1027 vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__nor2_4
XANTENNA__10107__B _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12145_ net255 net2480 net513 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__mux2_1
XANTENNA__09781__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09208__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16953_ clknet_leaf_151_wb_clk_i _02622_ _01182_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[926\]
+ sky130_fd_sc_hd__dfrtp_1
X_12076_ net239 net676 vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__and2_2
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ team_04_WB.MEM_SIZE_REG_REG\[27\] team_04_WB.MEM_SIZE_REG_REG\[26\] _06515_
+ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__or3_1
X_15904_ clknet_leaf_11_wb_clk_i _01581_ _00131_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16884_ clknet_leaf_2_wb_clk_i _02553_ _01113_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[857\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835_ clknet_leaf_88_wb_clk_i _01512_ _00062_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15766_ net1291 vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__inv_2
XANTENNA__11880__C _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12978_ net601 _07386_ net468 net314 net1675 vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a32o_1
XANTENNA__09123__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717_ net1149 vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11929_ net687 _07392_ _07394_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15697_ net1269 vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14648_ net1207 vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_70_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_28 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_39 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ net1259 vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16318_ clknet_leaf_158_wb_clk_i _01987_ _00547_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17298_ net1354 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13148__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16249_ clknet_leaf_154_wb_clk_i _01918_ _00478_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__B1 _07622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput135 net135 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__clkbuf_4
Xoutput146 net146 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput157 net157 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
Xoutput168 net168 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__clkbuf_4
XANTENNA_max_cap804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput179 net179 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10732__S net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07953_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net973 _03562_ vssd1 vssd1 vccd1
+ vccd1 _03564_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08202__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13856__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08958__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[10\] vssd1 vssd1
+ vccd1 vccd1 _03499_ sky130_fd_sc_hd__inv_2
XANTENNA__09822__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _05230_ _05231_ _05232_ _05233_ net834 net738 vssd1 vssd1 vccd1 vccd1 _05234_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12659__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13344__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ _05159_ _05164_ net775 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08505_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[311\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[279\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__mux2_1
X_09485_ _05092_ _05093_ _05094_ _05095_ net792 net802 vssd1 vssd1 vccd1 vccd1 _05096_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[952\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[920\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_77_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[377\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[345\]
+ net911 vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout322_X net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08444__Y _04055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09460__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08298_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[859\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13139__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09438__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ _05567_ _05641_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09763__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _05541_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\]
+ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10642__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout340 net341 vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout351 _07667_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
Xfanout362 _06253_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
X_13950_ _05467_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nor2_1
Xfanout373 net374 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
Xfanout384 _07674_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_8
Xfanout395 _07672_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_2
XANTENNA__09732__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ _07603_ net332 net384 net2203 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__a22o_1
X_13881_ _02910_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__nand2_1
XANTENNA__11873__A2 _07346_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__A net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ net1171 vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12832_ _07530_ net327 net392 net1748 vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08177__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15551_ net1270 vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__inv_2
XANTENNA__11625__A2 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12763_ _07490_ net334 net397 net1691 vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14502_ net1263 vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__inv_2
X_11714_ _06956_ _06957_ _06975_ _06976_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15482_ net1144 vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__inv_2
X_12694_ net2121 net406 net340 _07265_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17221_ net1427 _02831_ _01469_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_14433_ net1291 vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__inv_2
X_11645_ _07103_ _07133_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09677__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__B1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17152_ clknet_leaf_84_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[6\]
+ _01381_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xinput15 DAT_I[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ net1444 vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__clkbuf_1
Xinput26 DAT_I[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_154_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12050__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ net555 _07063_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__o21ai_1
Xinput37 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12317__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput48 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_16103_ clknet_leaf_24_wb_clk_i _01772_ _00332_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput59 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
X_13315_ net1084 team_04_WB.MEM_SIZE_REG_REG\[21\] vssd1 vssd1 vccd1 vccd1 _07741_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__14327__A1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17083_ clknet_leaf_43_wb_clk_i _00039_ _01312_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter_state
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net1095 net1054 vssd1 vssd1 vccd1
+ vccd1 _06090_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[27\] _03462_
+ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and2_1
XFILLER_0_126_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08006__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16034_ clknet_leaf_144_wb_clk_i _01703_ _00263_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_13246_ net92 net2663 net975 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__mux2_1
X_10458_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_90_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10349__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10389_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _05526_ vssd1
+ vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13177_ _07613_ net370 net290 net1644 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a22o_1
XANTENNA__12333__A _07374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09118__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ net212 net2482 net513 vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
X_12059_ net436 net676 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__nand2_4
X_16936_ clknet_leaf_114_wb_clk_i _02605_ _01165_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12620__X _07661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08957__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09601__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__B net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ clknet_leaf_124_wb_clk_i _02536_ _01096_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10788__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ clknet_leaf_88_wb_clk_i _01495_ _00045_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_16798_ clknet_leaf_116_wb_clk_i _02467_ _01027_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[771\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15749_ net1275 vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09270_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[841\]
+ net923 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__mux2_1
XANTENNA__09788__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_738 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08221_ _03828_ _03829_ _03830_ _03831_ net791 net812 vssd1 vssd1 vccd1 vccd1 _03832_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13611__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12577__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__A team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08152_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[188\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\]
+ net946 vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08083_ _03645_ _03693_ net663 vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__mux2_2
XANTENNA__12942__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_124_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_139_82 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08985_ _04592_ _04593_ _04594_ _04595_ net796 net803 vssd1 vssd1 vccd1 vccd1 _04596_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout484_A net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ net1079 net1028 net1024 vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__and3_1
XANTENNA__09823__Y _05434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12501__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_X net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout651_A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout749_A net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09606_ _05213_ _05214_ _05215_ _05216_ net793 net802 vssd1 vssd1 vccd1 vccd1 _05217_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08168__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09537_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[229\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\]
+ net956 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1181_X net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_A net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1279_X net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[742\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__inv_2
XANTENNA__10637__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _05006_ _05007_ _05008_ _05009_ net833 net738 vssd1 vssd1 vccd1 vccd1 _05010_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12568__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _06357_ _06445_ _06453_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08107__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09433__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12032__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__B2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ _06246_ _06615_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13780__A2 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10312_ _05583_ _05632_ net619 vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__a21o_1
XANTENNA__11791__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ _07532_ net367 net298 net1923 vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__a22o_1
XANTENNA__09727__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14080_ net1467 _06106_ net1032 vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__mux2_1
X_11292_ net463 _06764_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_105_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10243_ _05538_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nor2_1
X_13031_ _07492_ net368 net306 net1596 vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__a22o_1
XANTENNA__13532__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input45_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1102 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\] vssd1
+ vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
X_10174_ _05543_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__nand2b_1
Xfanout1113 net1114 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__buf_4
Xfanout1124 net1127 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__buf_4
Xfanout1135 net1157 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_2
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_4
XANTENNA__08777__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14982_ net1103 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__inv_2
XANTENNA__12099__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1157 net1158 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_2
XANTENNA__12440__X _07641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1168 net1169 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__clkbuf_4
X_16721_ clknet_leaf_172_wb_clk_i _02390_ _00950_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\]
+ sky130_fd_sc_hd__dfrtp_1
X_13933_ _03094_ net1040 _03298_ net1071 net131 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a32o_1
XANTENNA__08398__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08172__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16652_ clknet_leaf_111_wb_clk_i _02321_ _00881_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\]
+ sky130_fd_sc_hd__dfrtp_1
X_13864_ _02886_ _02895_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__or3_1
X_15603_ net1232 vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ net261 net2303 net324 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__mux2_1
XANTENNA__09347__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output201_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16583_ clknet_leaf_21_wb_clk_i _02252_ _00812_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\]
+ sky130_fd_sc_hd__dfrtp_1
X_13795_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] _05896_ net1100
+ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13712__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10806__B1 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15534_ net1203 vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__inv_2
X_12746_ _07471_ net328 net400 net2277 vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__a22o_1
XANTENNA__12271__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13633__A2_N net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09401__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10282__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10547__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15465_ net1135 vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12677_ net250 net2618 net478 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ net1410 _02814_ _01435_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_13_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416_ net1283 vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11628_ team_04_WB.MEM_SIZE_REG_REG\[1\] _07116_ vssd1 vssd1 vccd1 vccd1 _07117_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15396_ net1183 vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__inv_2
XANTENNA__12047__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17135_ clknet_leaf_82_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[0\]
+ _01364_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ net1191 vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ net565 _07043_ _07044_ net570 vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__a31o_1
XANTENNA__11782__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\] vssd1 vssd1
+ vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold618 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\] vssd1 vssd1
+ vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ clknet_leaf_48_wb_clk_i _00013_ _01295_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold629 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\] vssd1 vssd1
+ vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14278_ _03452_ net819 _03451_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__and3b_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16017_ clknet_leaf_52_wb_clk_i _01693_ _00246_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_59_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13229_ net72 team_04_WB.MEM_SIZE_REG_REG\[12\] net984 vssd1 vssd1 vccd1 vccd1 _01674_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11534__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12731__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6__f_wb_clk_i clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08770_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[690\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__mux2_1
XANTENNA__08687__S net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16919_ clknet_leaf_173_wb_clk_i _02588_ _01148_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[892\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13039__A1 _07500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12937__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09322_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08716__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ _04846_ _04852_ _04863_ net716 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a22o_4
XFILLER_0_157_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout232_A _07420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12238__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08204_ _03811_ _03812_ _03813_ _03814_ net791 net812 vssd1 vssd1 vccd1 vccd1 _03815_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09184_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12014__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_170_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08135_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__mux2_1
XANTENNA__12672__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11773__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12970__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12404__C net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12722__B1 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__X _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15284__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08597__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__mux2_1
XANTENNA__09282__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nand2_1
XANTENNA__08169__Y _03780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10930_ net588 _06399_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_92_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_169_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09329__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ _06348_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_21_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ _07569_ net484 net413 net2091 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__a22o_1
XANTENNA__12789__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08048__D net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13580_ _06900_ net272 net710 vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__a21o_1
XANTENNA__12253__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10792_ net586 _06207_ _06225_ _06276_ net287 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__o311a_1
XFILLER_0_151_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09221__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12531_ net2217 net247 net420 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15250_ net1246 vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_12462_ net522 net603 _07463_ net429 net1629 vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a32o_1
XANTENNA__09406__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__inv_2
X_11413_ _06507_ _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_590 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ net1199 vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ net521 _07247_ net603 net432 net1841 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14132_ team_04_WB.MEM_SIZE_REG_REG\[31\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[31\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__o221a_1
XFILLER_0_151_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11764__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12961__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _06246_ _06831_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14063_ net2 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1
+ vccd1 vccd1 _01523_ sky130_fd_sc_hd__o22a_1
X_11275_ _06468_ _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12713__B1 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_148_Right_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13014_ net608 _07474_ net472 net312 net1723 vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a32o_1
X_10226_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _05539_ vssd1
+ vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__xor2_1
XANTENNA__08393__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _05679_ _05767_ _05677_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\] vssd1 vssd1 vccd1
+ vccd1 net1441 sky130_fd_sc_hd__dlygate4sd3_1
X_10088_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _04559_ vssd1
+ vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__nand2_1
X_14965_ net1201 vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13916_ _03098_ _03142_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__or2_1
X_16704_ clknet_leaf_139_wb_clk_i _02373_ _00933_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14896_ net1173 vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__inv_2
XANTENNA__09893__B1 _04166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16635_ clknet_leaf_100_wb_clk_i _02304_ _00864_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[608\]
+ sky130_fd_sc_hd__dfrtp_1
X_13847_ net992 _03235_ _03237_ net990 vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_18_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16566_ clknet_leaf_15_wb_clk_i _02235_ _00795_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\]
+ sky130_fd_sc_hd__dfrtp_1
X_13778_ team_04_WB.ADDR_START_VAL_REG\[18\] _03167_ vssd1 vssd1 vccd1 vccd1 _03169_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09131__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_wb_clk_i_X clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15517_ net1153 vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12729_ _07454_ net333 net401 net2289 vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
X_16497_ clknet_leaf_179_wb_clk_i _02166_ _00726_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15448_ net1221 vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15379_ net1246 vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11755__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17118_ clknet_leaf_65_wb_clk_i _02753_ _01347_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold404 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\] vssd1 vssd1
+ vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08620__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold415 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\] vssd1 vssd1
+ vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\] vssd1 vssd1
+ vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold437 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\] vssd1 vssd1
+ vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold448 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[212\] vssd1 vssd1
+ vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__nand2_1
X_17049_ clknet_leaf_178_wb_clk_i _02718_ _01278_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold459 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\] vssd1 vssd1
+ vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12704__B1 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout906 net907 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout917 net920 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__clkbuf_4
X_09871_ _05032_ _05057_ _05084_ _05030_ _05004_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__o32a_1
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_2
XANTENNA__12180__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12080__X _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\] vssd1 vssd1
+ vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\] vssd1 vssd1
+ vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[158\] vssd1 vssd1
+ vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09306__S net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1137 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\] vssd1 vssd1
+ vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ _04360_ _04361_ _04362_ _04363_ net787 net810 vssd1 vssd1 vccd1 vccd1 _04364_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__17092__Q team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1148 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\] vssd1 vssd1
+ vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\] vssd1 vssd1
+ vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12240__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08684_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__B1 _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12667__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout447_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__Y _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12235__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_172_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09041__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _04912_ _04913_ _04914_ _04915_ net826 net742 vssd1 vssd1 vccd1 vccd1 _04916_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11994__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ _04772_ _04777_ net772 vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12943__A0 _07374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[382\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[350\]
+ net851 vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[45\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[13\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout983_A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08049_ net1078 net1030 net1026 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\]
+ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__o31a_1
Xhold960 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[976\] vssd1 vssd1
+ vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14911__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold971 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\] vssd1 vssd1
+ vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[785\] vssd1 vssd1
+ vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ _04328_ net549 vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nand2_1
Xhold993 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\] vssd1 vssd1
+ vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ net627 _04948_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10503__X _06073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09216__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08120__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ net1217 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11962_ _03631_ _05988_ net696 _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__a211o_1
XANTENNA__13671__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__B2 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10913_ net570 net657 _06269_ _06401_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__o211a_1
XFILLER_0_169_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14681_ net1237 vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__inv_2
XANTENNA__14358__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07364_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_80_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16420_ clknet_leaf_165_wb_clk_i _02089_ _00649_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13632_ _07076_ net271 _07687_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__a22o_1
X_17333__1389 vssd1 vssd1 vccd1 vccd1 _17333__1389/HI net1389 sky130_fd_sc_hd__conb_1
X_10844_ _04029_ _06305_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16351_ clknet_leaf_155_wb_clk_i _02020_ _00580_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[324\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08525__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ net998 _02953_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__nand2_1
X_10775_ _03721_ net550 vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11985__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ net1104 vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__inv_2
X_12514_ _07511_ net490 net426 net1598 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08790__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16282_ clknet_leaf_37_wb_clk_i _01951_ _00511_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\]
+ sky130_fd_sc_hd__dfrtp_1
X_13494_ _02876_ _02880_ _02883_ team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1
+ vccd1 _02885_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output199_A net199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__B1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15233_ net1169 vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__inv_2
X_12445_ net2452 net430 _07643_ net523 vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12934__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15164_ net1148 vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12376_ _07356_ net2459 net497 vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__mux2_1
X_17243__1405 vssd1 vssd1 vccd1 vccd1 net1405 _17243__1405/LO sky130_fd_sc_hd__conb_1
XANTENNA__12325__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ team_04_WB.MEM_SIZE_REG_REG\[14\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[14\]
+ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__a22o_1
X_11327_ net753 _06786_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__and3_2
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10126__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15095_ net1231 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14046_ net10 net1063 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1
+ vccd1 vccd1 _01540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ _06745_ _06746_ net567 vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12162__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10209_ _05541_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11189_ net582 _06677_ net288 vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09126__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15997_ clknet_leaf_69_wb_clk_i _01673_ _00226_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12060__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13111__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14948_ net1189 vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12465__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14879_ net1265 vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ clknet_leaf_163_wb_clk_i _02287_ _00847_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12059__Y _07484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16549_ clknet_leaf_185_wb_clk_i _02218_ _00778_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13965__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__B1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11976__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11440__A3 _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13178__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09021_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[878\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[846\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12925__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold201 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[191\] vssd1 vssd1
+ vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold212 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\] vssd1 vssd1
+ vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[615\] vssd1 vssd1
+ vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14127__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10400__A1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold234 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[371\] vssd1 vssd1
+ vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12950__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[618\] vssd1 vssd1
+ vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold256 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[686\] vssd1 vssd1
+ vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold267 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[367\] vssd1 vssd1
+ vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold278 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\] vssd1 vssd1
+ vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\]
+ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_113_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09825__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout703 _03642_ vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
Xhold289 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\] vssd1 vssd1
+ vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 net715 vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout397_A _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 net726 vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13347__A team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout736 net740 vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout747 net749 vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
X_09854_ _05460_ net659 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__or2_1
Xfanout758 _03613_ vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07990__D net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1104_A net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 _03569_ vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__buf_4
XANTENNA__11900__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__S net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[273\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09785_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\]
+ net961 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout564_A net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
XANTENNA__08204__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__B1 _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout731_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12208__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09085__A1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1261_X net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10560_ team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] net1095 net1051 vssd1 vssd1 vccd1
+ vccd1 _06112_ sky130_fd_sc_hd__and3_1
XFILLER_0_107_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13169__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13708__A2 _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[938\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10491_ _06028_ _06037_ _06049_ _06051_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__and4_1
XANTENNA__12426__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12916__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12230_ net213 net674 vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ net211 net648 vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11112_ net545 _06531_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12092_ net258 net678 vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__and2_1
Xhold790 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\] vssd1 vssd1
+ vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15920_ clknet_leaf_73_wb_clk_i _01597_ _00147_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11043_ net645 net571 vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__nor2_2
XANTENNA__12161__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12695__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ clknet_leaf_86_wb_clk_i _01528_ _00078_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_14802_ net1244 vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__inv_2
X_15782_ net1287 vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__inv_2
XANTENNA__12447__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _07645_ net470 net311 net2144 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10112__C _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ net1210 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11945_ net653 net234 vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14664_ net1117 vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__inv_2
X_11876_ net656 net259 vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_60_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16403_ clknet_leaf_182_wb_clk_i _02072_ _00632_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[376\]
+ sky130_fd_sc_hd__dfrtp_1
X_13615_ _07785_ _07800_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10827_ _03861_ _06310_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__xnor2_1
X_14595_ net1176 vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__inv_2
XANTENNA__14816__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11958__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ clknet_leaf_26_wb_clk_i _02003_ _00563_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[307\]
+ sky130_fd_sc_hd__dfrtp_1
X_13546_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\] net1043 _02936_
+ net1081 vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_45_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10758_ net568 _06207_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__or2_2
XFILLER_0_54_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08814__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16265_ clknet_leaf_121_wb_clk_i _01934_ _00494_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[28\] net1043 _02867_
+ net1092 vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10555__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10689_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[3\] net711 _06180_
+ net2273 vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15216_ net1163 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__inv_2
XANTENNA__12907__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ net654 net608 net224 vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__and3_1
X_16196_ clknet_leaf_168_wb_clk_i _01865_ _00425_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[169\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12055__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13580__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15147_ net1167 vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12359_ _06194_ _07249_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__or2_4
XFILLER_0_121_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14124__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15078_ net1103 vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_68 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029_ net1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03351_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_71_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09000__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08985__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[805\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_160_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08695__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08521_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__mux2_1
XANTENNA__08737__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_149_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_149_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08452_ net720 _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13938__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08383_ _03990_ _03991_ _03992_ _03993_ net783 net805 vssd1 vssd1 vccd1 vccd1 _03994_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12945__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13630__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08283__X _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12610__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10621__A1 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_115_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_167_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12680__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14461__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_105_wb_clk_i_A clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14115__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332__1388 vssd1 vssd1 vccd1 vccd1 _17332__1388/HI net1388 sky130_fd_sc_hd__conb_1
XFILLER_0_111_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout500 _07591_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_4
XANTENNA_fanout681_A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout779_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net512 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__buf_6
X_09906_ _05439_ _05509_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nand2_1
Xfanout522 _06197_ vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_4
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
XFILLER_0_158_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08425__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13874__B2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 net556 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__buf_2
X_09837_ _04784_ _05443_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__nand2_1
Xfanout577 net578 vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11885__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout588 _05110_ vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_2
Xfanout599 _03309_ vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_4
XANTENNA__12429__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _05336_ net551 vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08719_ _03640_ _03644_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__and2_2
XFILLER_0_69_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ net664 _05307_ _05308_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08502__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11730_ _06816_ _06817_ _06935_ _06955_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_166_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11661_ net463 _07141_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__o21ai_2
XANTENNA__09058__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14051__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_13400_ net1085 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 _07826_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_25_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11612__X _07101_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ net53 net52 net55 net54 vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_25_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14380_ net1497 vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12601__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11592_ _05312_ _06248_ _06253_ _05311_ _07080_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_144_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _07753_ _07755_ _07756_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[19\]
+ _06100_ net1047 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11060__A _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16050_ clknet_leaf_7_wb_clk_i _01719_ _00279_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input75_A wbs_dat_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ net74 team_04_WB.ADDR_START_VAL_REG\[14\] net976 vssd1 vssd1 vccd1 vccd1
+ _01644_ sky130_fd_sc_hd__mux2_1
X_10474_ _06037_ _06049_ _06051_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_40_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08569__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15001_ net1239 vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__inv_2
X_12213_ net224 net649 vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__and2_1
XANTENNA__11995__A net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ net1028 net1027 vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10107__C _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14106__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ net256 net2504 net514 vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16952_ clknet_leaf_148_wb_clk_i _02621_ _01181_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[925\]
+ sky130_fd_sc_hd__dfrtp_1
X_12075_ net2237 net352 _07492_ net440 vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a22o_1
X_11026_ team_04_WB.MEM_SIZE_REG_REG\[25\] _06514_ vssd1 vssd1 vccd1 vccd1 _06515_
+ sky130_fd_sc_hd__or2_1
X_15903_ clknet_leaf_11_wb_clk_i _01580_ _00130_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__dfrtp_1
XANTENNA__10679__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16883_ clknet_leaf_181_wb_clk_i _02552_ _01112_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13715__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15834_ clknet_leaf_89_wb_clk_i _01511_ _00061_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09912__B _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15765_ net1291 vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
X_12977_ net601 _07381_ net469 net314 net1568 vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13093__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_183_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11928_ net759 _05952_ net695 _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_47_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14716_ net1126 vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15696_ net1268 vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12840__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_72_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14647_ net1223 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11859_ net1910 net527 net447 _07334_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a22o_1
XANTENNA__14546__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14042__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_18 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578_ net1259 vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_29 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10793__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13529_ team_04_WB.ADDR_START_VAL_REG\[22\] _02918_ vssd1 vssd1 vccd1 vccd1 _02920_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16317_ clknet_leaf_129_wb_clk_i _01986_ _00546_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17297_ net1353 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XFILLER_0_166_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16248_ clknet_leaf_153_wb_clk_i _01917_ _00477_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__clkbuf_4
X_16179_ clknet_leaf_185_wb_clk_i _01848_ _00408_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput125 net125 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08655__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput136 net136 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
Xoutput147 net147 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_81_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput158 net158 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
Xoutput169 net169 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__13609__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07952_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net973 _03562_ vssd1 vssd1 vccd1
+ vccd1 _03563_ sky130_fd_sc_hd__o21a_1
XANTENNA__08958__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11867__B1 net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07883_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\] vssd1 vssd1
+ vccd1 vccd1 _03498_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08732__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[35\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__mux2_1
XANTENNA__08719__A _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09314__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _05160_ _05161_ _05162_ _05163_ net793 net813 vssd1 vssd1 vccd1 vccd1 _05164_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_108_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout262_A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08504_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[343\]
+ net845 vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__mux2_1
XANTENNA__11095__A1 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__mux2_1
XANTENNA__12831__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__mux2_1
XANTENNA__12675__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14033__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout527_A _06195_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1269_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ net642 _03974_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_163_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13792__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09460__A1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1057_X net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout896_A net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ net622 _05797_ _05796_ net281 vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13847__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_4
Xfanout341 net351 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 net353 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_6
XANTENNA__11039__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout363 net365 vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09071__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 _07674_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_4
X_12900_ _07602_ net326 net384 net1892 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a22o_1
Xfanout396 _07670_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_6
X_13880_ _02921_ _02932_ _03260_ _02919_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a31o_1
XANTENNA__09224__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ _07529_ net329 net392 net1766 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a22o_1
XANTENNA__11055__A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15550_ net1216 vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__inv_2
X_12762_ _07489_ net333 net397 net1944 vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ net1285 vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11713_ _06732_ _06818_ _06881_ _06841_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15481_ net1251 vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__inv_2
X_12693_ net2257 net406 net340 _07259_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17220_ net1426 _02830_ _01467_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[20\]
+ sky130_fd_sc_hd__dfrtp_2
X_14432_ net1277 vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__inv_2
X_11644_ team_04_WB.MEM_SIZE_REG_REG\[3\] team_04_WB.MEM_SIZE_REG_REG\[2\] vssd1 vssd1
+ vccd1 vccd1 _07133_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_42_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17151_ clknet_leaf_84_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[5\]
+ _01380_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_3_5_0_wb_clk_i_X clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ net1554 vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11575_ net564 _06985_ net577 vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o21a_1
Xinput16 DAT_I[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_17239__1300 vssd1 vssd1 vccd1 vccd1 _17239__1300/HI net1300 sky130_fd_sc_hd__conb_1
Xinput27 DAT_I[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16102_ clknet_leaf_19_wb_clk_i _01771_ _00331_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput38 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_1
X_13314_ net1083 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 _07740_
+ sky130_fd_sc_hd__nand2_1
Xinput49 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
X_10526_ _06089_ net1614 net1022 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
X_17082_ clknet_leaf_45_wb_clk_i net2641 _01311_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14294_ _03462_ net818 _03461_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__and3b_1
XANTENNA_output181_A net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__B _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ clknet_leaf_136_wb_clk_i _01702_ _00262_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12338__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ net93 team_04_WB.ADDR_START_VAL_REG\[31\] net976 vssd1 vssd1 vccd1 vccd1
+ _01661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_131_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15197__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ _06034_ _06035_ _06030_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_131_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08006__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13176_ _07612_ net370 net290 net1655 vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__a22o_1
XANTENNA__08303__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ net623 _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__nor2_1
XANTENNA__12333__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _07246_ net2502 net512 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_16935_ clknet_leaf_165_wb_clk_i _02604_ _01164_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\]
+ sky130_fd_sc_hd__dfrtp_1
X_12058_ _04783_ _05280_ net822 vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__or3_1
XANTENNA__11313__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net464 _06496_ _06497_ _06281_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a31o_2
XFILLER_0_74_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16866_ clknet_leaf_146_wb_clk_i _02535_ _01095_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10788__B _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15817_ clknet_leaf_89_wb_clk_i _01494_ _00044_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_16797_ clknet_leaf_126_wb_clk_i _02466_ _01026_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ net1275 vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__inv_2
XANTENNA__08973__S net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15679_ net1281 vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331__1387 vssd1 vssd1 vccd1 vccd1 _17331__1387/HI net1387 sky130_fd_sc_hd__conb_1
XFILLER_0_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08220_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[701\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[669\]
+ net950 vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08151_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[252\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\]
+ net946 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08082_ _03672_ _03681_ _03692_ net717 vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__a22o_2
XFILLER_0_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08280__Y _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08213__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08984_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[46\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_94 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1017_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ net1054 _03543_ _03544_ _03535_ _03537_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__o221ai_2
Xclkbuf_leaf_164_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_164_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout477_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1059 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09605_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[547\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09536_ _05143_ _05144_ _05145_ _05146_ net793 net813 vssd1 vssd1 vccd1 vccd1 _05147_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout811_A _03550_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout909_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11162__X _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08418_ _04004_ _04028_ net663 vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__mux2_2
XFILLER_0_47_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[295\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[263\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_478 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ net722 _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__or2_1
XANTENNA__09433__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Left_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11240__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11360_ _06607_ _06619_ net569 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13780__A3 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11749__S net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] net1075 _05903_
+ _05905_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__o22a_1
XANTENNA__13089__X _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09727__B net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08619__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11291_ net286 _06775_ _06779_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__or3_2
XANTENNA__12434__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11528__C1 _07016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09219__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ _07491_ net367 net306 net2018 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__a22o_1
X_10242_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[21\] _05537_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10200__C1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10173_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[29\] _05542_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\]
+ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__a21o_1
Xfanout1103 net1115 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__buf_4
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1114 net1115 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
Xfanout1125 net1127 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__buf_2
Xfanout1136 net1138 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__buf_4
XANTENNA_input38_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1147 net1156 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
X_14981_ net1113 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__inv_2
Xfanout1158 net1194 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_137_Left_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1169 net1187 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16720_ clknet_leaf_191_wb_clk_i _02389_ _00949_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[693\]
+ sky130_fd_sc_hd__dfrtp_1
X_13932_ _03018_ _03093_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__nand2_1
XANTENNA__08172__A1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ _03222_ _03223_ _02897_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__o21a_1
X_16651_ clknet_leaf_31_wb_clk_i _02320_ _00880_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13048__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ net1245 vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__inv_2
X_12814_ net249 net2406 net325 vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__mux2_1
XANTENNA__09347__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] net1044 _03184_
+ net1081 vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o22a_1
X_16582_ clknet_leaf_22_wb_clk_i _02251_ _00811_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15533_ net1144 vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__inv_2
X_12745_ _07470_ net333 net401 net2398 vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09672__A1 _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11072__X _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15464_ net1117 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__inv_2
X_12676_ net251 net2138 net475 vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_146_Left_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ net1409 _02813_ _01433_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_133_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ net1267 vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11627_ net754 _07115_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15395_ net1182 vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08858__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17134_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[1\]
+ _01363_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_14346_ net1191 vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ net532 _07046_ _07045_ net556 vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11782__A2 _05800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\] vssd1 vssd1
+ vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ clknet_leaf_49_wb_clk_i _00012_ _01294_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10509_ team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] net1097 net1053 vssd1 vssd1 vccd1
+ vccd1 _06078_ sky130_fd_sc_hd__and3_1
X_14277_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\]
+ _03448_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and3_1
Xhold619 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\] vssd1 vssd1
+ vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ _06442_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__nand2_1
X_16016_ clknet_leaf_52_wb_clk_i _01692_ _00245_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09188__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ net73 team_04_WB.MEM_SIZE_REG_REG\[13\] net983 vssd1 vssd1 vccd1 vccd1 _01675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08033__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13159_ _07595_ net377 net292 net1926 vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10742__A0 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_155_Left_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16918_ clknet_leaf_11_wb_clk_i _02587_ _01147_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12495__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
X_16849_ clknet_leaf_180_wb_clk_i _02518_ _01078_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13039__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09799__S net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_157_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07901__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\]
+ net960 vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ _04857_ _04862_ net720 vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08208__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12238__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[413\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12953__S net321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_170_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08134_ _03741_ _03742_ _03743_ _03744_ net831 net737 vssd1 vssd1 vccd1 vccd1 _03745_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12970__A1 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\]
+ net865 vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__mux2_1
XANTENNA__12254__A net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09039__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09274__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout594_A _04112_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10733__A0 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout761_A _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout382_X net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__inv_2
XANTENNA__12486__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08898_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\]
+ net872 vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout647_X net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ _04218_ _06347_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nand2_1
XANTENNA__09329__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _05126_ _05127_ _05128_ _05129_ net831 net747 vssd1 vssd1 vccd1 vccd1 _05130_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _05464_ _06277_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12530_ net2196 net240 net421 vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08118__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12461_ net522 net604 _07462_ net429 net1667 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a32o_1
XANTENNA__09406__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1090
+ net1089 vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__and3_1
X_11412_ team_04_WB.MEM_SIZE_REG_REG\[13\] _06506_ vssd1 vssd1 vccd1 vccd1 _06901_
+ sky130_fd_sc_hd__nand2_1
X_15180_ net1121 vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__inv_2
XANTENNA__09738__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ net699 _06183_ _06198_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__or3_4
XANTENNA__11987__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14131_ team_04_WB.MEM_SIZE_REG_REG\[30\] net988 net981 team_04_WB.ADDR_START_VAL_REG\[30\]
+ net1005 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__o221a_1
XANTENNA__11764__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ net562 _05475_ _06240_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__and3_1
XFILLER_0_105_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ net13 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1 vssd1
+ vccd1 vccd1 _01524_ sky130_fd_sc_hd__a22o_1
X_11274_ _04501_ _06356_ _06454_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_37_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13013_ net611 _07473_ net474 net313 net2340 vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a32o_1
XANTENNA__13910__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ _05648_ net621 _05826_ _05828_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11921__C1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17330__1386 vssd1 vssd1 vccd1 vccd1 _17330__1386/HI net1386 sky130_fd_sc_hd__conb_1
X_10156_ _05681_ _05765_ _05680_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a21boi_1
XANTENNA__09017__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output144_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 net139 vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__inv_2
X_14964_ net1235 vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ clknet_leaf_157_wb_clk_i _02372_ _00932_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[676\]
+ sky130_fd_sc_hd__dfrtp_1
X_13915_ _03243_ _03286_ net1696 net1071 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_50_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__A1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14895_ net1140 vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__inv_2
XANTENNA__11942__S _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16634_ clknet_leaf_38_wb_clk_i _02303_ _00863_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\]
+ sky130_fd_sc_hd__dfrtp_1
X_13846_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] _05544_ net1100
+ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09412__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ team_04_WB.ADDR_START_VAL_REG\[18\] _03167_ vssd1 vssd1 vccd1 vccd1 _03168_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10558__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16565_ clknet_leaf_15_wb_clk_i _02234_ _00794_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_168_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10989_ _06477_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__inv_2
XANTENNA__12339__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10255__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15516_ net1145 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
X_12728_ _07453_ net331 net400 net2132 vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16496_ clknet_leaf_192_wb_clk_i _02165_ _00725_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[469\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15447_ net1230 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__inv_2
X_12659_ net227 net2510 net476 vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15378_ net1247 vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07959__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11755__A2 _07242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17117_ clknet_leaf_104_wb_clk_i _02752_ _01346_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_14329_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[3\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[2\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[0\] net1090
+ net1089 vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__mux4_1
XANTENNA__10293__S net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\] vssd1 vssd1
+ vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold416 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[227\] vssd1 vssd1
+ vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold427 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\] vssd1 vssd1
+ vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[114\] vssd1 vssd1
+ vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[223\] vssd1 vssd1
+ vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
X_17048_ clknet_leaf_150_wb_clk_i _02717_ _01277_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13901__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout907 net910 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__clkbuf_4
X_09870_ _05478_ _05480_ _05195_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a21bo_1
Xfanout918 net920 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08698__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout929 net941 vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12180__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08821_ net776 _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_146_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\] vssd1 vssd1
+ vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1116 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\] vssd1 vssd1
+ vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
Xhold1127 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[153\] vssd1 vssd1
+ vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10322__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1138 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\] vssd1 vssd1
+ vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1149 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[407\] vssd1 vssd1
+ vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08683_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[565\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
XANTENNA__12948__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__A2 net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09322__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11979__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[681\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[649\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_172_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12640__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11994__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09235_ net720 _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12683__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14464__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1251_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09166_ _04773_ _04774_ _04775_ _04776_ net789 net800 vssd1 vssd1 vccd1 vccd1 _04777_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08117_ net752 _03727_ _03726_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_82_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_1__f_wb_clk_i_A clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08048_ _03510_ net1078 net1030 net1026 vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or4_4
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold950 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\] vssd1 vssd1
+ vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout976_A net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[459\] vssd1 vssd1
+ vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\] vssd1 vssd1
+ vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold983 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\] vssd1 vssd1
+ vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[725\] vssd1 vssd1
+ vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _05598_ _05620_ _05597_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08401__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _05276_ _05282_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09580__X _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ net756 _05989_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ _03032_ _03089_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__nor2_1
X_10912_ net576 net659 _06226_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or3_1
X_14680_ net1203 vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__inv_2
XANTENNA__08196__X _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ net2126 net529 net458 _07363_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a22o_1
XANTENNA__08637__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09232__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13631_ _03540_ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10843_ _06328_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__and2_1
XANTENNA__10378__S net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13562_ net990 _02952_ _02950_ net995 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_149_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10237__A2 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16350_ clknet_leaf_115_wb_clk_i _02019_ _00579_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[323\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ net538 _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ _07510_ net490 net426 net1846 vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
X_15301_ net1108 vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16281_ clknet_leaf_154_wb_clk_i _01950_ _00510_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ team_04_WB.ADDR_START_VAL_REG\[27\] _02876_ _02880_ _02883_ vssd1 vssd1 vccd1
+ vccd1 _02884_ sky130_fd_sc_hd__and4_1
XFILLER_0_137_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ net607 net214 net682 vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15232_ net1211 vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ net1113 vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12375_ net259 net2642 net496 vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ team_04_WB.MEM_SIZE_REG_REG\[13\] net986 net979 team_04_WB.ADDR_START_VAL_REG\[13\]
+ net1003 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__o221a_1
X_11326_ net286 _06811_ _06814_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15094_ net1228 vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__inv_2
X_14045_ net11 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1
+ vccd1 vccd1 _01541_ sky130_fd_sc_hd__a22o_1
X_11257_ _06576_ _06582_ net562 vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__mux2_1
XANTENNA__14313__S net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12698__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10208_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\] _05540_ vssd1
+ vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__nor2_1
XANTENNA__12162__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08311__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17193__Q team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ net566 _06666_ _06536_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__o21a_1
XANTENNA__12341__B net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10139_ _05713_ _05749_ _05711_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15996_ clknet_leaf_69_wb_clk_i _01672_ _00225_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_14947_ net1170 vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12870__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14878_ net1239 vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__inv_2
XANTENNA__09142__S net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16617_ clknet_leaf_123_wb_clk_i _02286_ _00846_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\]
+ sky130_fd_sc_hd__dfrtp_1
X_13829_ team_04_WB.ADDR_START_VAL_REG\[24\] _03218_ vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10228__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12622__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16548_ clknet_leaf_171_wb_clk_i _02217_ _00777_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08981__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13965__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11976__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16479_ clknet_leaf_160_wb_clk_i _02148_ _00708_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13178__A1 _07614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09020_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[910\]
+ net901 vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold202 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\] vssd1 vssd1
+ vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold213 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\] vssd1 vssd1
+ vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14127__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__X _05276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\] vssd1 vssd1
+ vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold235 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\] vssd1 vssd1
+ vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold246 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\] vssd1 vssd1
+ vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_698 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold257 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\] vssd1 vssd1
+ vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold268 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\] vssd1 vssd1
+ vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[14\] _05532_ vssd1
+ vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and2_1
Xhold279 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[247\] vssd1 vssd1
+ vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_2
Xfanout715 _03675_ vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__buf_4
Xfanout726 _03668_ vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_165_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout737 net739 vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__clkbuf_8
X_09853_ _05460_ net658 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_165_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 net749 vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08804_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[369\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\]
+ net971 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__mux2_1
X_09784_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\]
+ net961 vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09841__A _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
XANTENNA__08204__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12678__S net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
XANTENNA__12861__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09052__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08597_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[788\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout345_X net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08744__X _04355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12613__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11967__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_134_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_X net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1254_X net1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13169__A1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09218_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[970\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10490_ _06047_ _06052_ _06064_ _06065_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__a31o_1
XANTENNA__13708__A3 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12426__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09149_ _04756_ _04757_ _04758_ _04759_ net784 net800 vssd1 vssd1 vccd1 vccd1 _04760_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_20_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14118__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ net701 _06194_ net650 vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11111_ net530 _06261_ _06264_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_9_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12091_ net2292 net353 _07500_ net446 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a22o_1
Xhold780 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\] vssd1 vssd1
+ vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12442__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold791 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\] vssd1 vssd1
+ vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ net645 net535 vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nor2_1
XANTENNA__08131__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12161__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ clknet_leaf_86_wb_clk_i _01527_ _00077_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_110_Left_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input20_A DAT_I[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ net1270 vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__inv_2
X_15781_ net1192 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__inv_2
X_12993_ _07644_ net473 net312 net2268 vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__a22o_1
XANTENNA__10897__A _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14732_ net1121 vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
X_11944_ net695 _07038_ _07407_ net616 vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__a211oi_2
XANTENNA_clkbuf_leaf_173_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12852__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875_ net613 _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__and3_2
X_14663_ net1134 vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__inv_2
X_16402_ clknet_leaf_9_wb_clk_i _02071_ _00631_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[375\]
+ sky130_fd_sc_hd__dfrtp_1
X_13614_ _02999_ _03002_ _03004_ team_04_WB.ADDR_START_VAL_REG\[7\] vssd1 vssd1 vccd1
+ vccd1 _03005_ sky130_fd_sc_hd__a31o_1
X_10826_ _06313_ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__nor2_1
XANTENNA__11407__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12604__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ net1184 vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__inv_2
XANTENNA__11958__A2 _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13720__B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ clknet_leaf_44_wb_clk_i _02002_ _00562_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\]
+ sky130_fd_sc_hd__dfrtp_1
X_13545_ _07840_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10757_ net569 _06207_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_45_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13212__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _07870_ _02866_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__nand2b_1
X_16264_ clknet_leaf_113_wb_clk_i _01933_ _00493_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[4\] net711 _06180_
+ net1701 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
XANTENNA__09459__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15215_ net1196 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__inv_2
X_12427_ net2003 net434 _07634_ net524 vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16195_ clknet_leaf_116_wb_clk_i _01864_ _00424_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14832__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14109__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__C net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12358_ net2208 net502 _07623_ net460 vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a22o_1
X_15146_ net1111 vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _06795_ _06797_ net560 vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__mux2_1
X_15077_ net1111 vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ net2585 net505 _07587_ net455 vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
X_14028_ net1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03350_ sky130_fd_sc_hd__and2_1
XANTENNA__09137__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0__f_wb_clk_i_X clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13883__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08976__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08829__X _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_160_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13096__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_160_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15979_ clknet_leaf_43_wb_clk_i _01655_ _00208_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08520_ _04127_ _04128_ _04129_ _04130_ net824 net733 vssd1 vssd1 vccd1 vccd1 _04131_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12843__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08451_ _04058_ _04059_ _04060_ _04061_ net825 net742 vssd1 vssd1 vccd1 vccd1 _04062_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08382_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[921\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_189_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_189_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09600__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_118_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_144_943 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12246__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[366\] net899 _03662_
+ _04613_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o211a_1
XFILLER_0_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10047__A net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout305_A _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_114 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08122__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_167_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12262__A net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout501 net502 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_8
X_09905_ _05514_ _05515_ _03866_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__o21ai_4
Xfanout512 net514 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_6
Xfanout523 net525 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_4
Xfanout534 _05435_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08425__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout674_A _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_X net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _05377_ vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
Xfanout556 _05310_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__buf_2
XANTENNA__10688__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 net568 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
X_09836_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08886__S net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout578 _05250_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_2
Xfanout589 _05003_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13087__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ net664 _05375_ _05340_ _05336_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__a211o_1
XANTENNA__08189__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08718_ net765 _04321_ _04327_ _04315_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__a31o_2
XANTENNA__11637__A1 _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ net664 _05307_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08649_ _04256_ _04257_ _04258_ _04259_ net783 net800 vssd1 vssd1 vccd1 vccd1 _04260_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _05473_ _07144_ _07147_ _07148_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09689__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09510__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ _06147_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11496__S0 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ net625 net555 _06257_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__and3b_1
XFILLER_0_147_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ net1086 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 _07756_
+ sky130_fd_sc_hd__nor2_1
X_10542_ team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] net1095 net1051 vssd1 vssd1 vccd1
+ vccd1 _06100_ sky130_fd_sc_hd__and3_1
XANTENNA__08126__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13261_ net75 team_04_WB.ADDR_START_VAL_REG\[15\] net975 vssd1 vssd1 vccd1 vccd1
+ _01645_ sky130_fd_sc_hd__mux2_1
X_10473_ _06050_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__and2_1
XANTENNA__13011__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__X _07669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__Y _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08569__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ net2261 net509 _07547_ net454 vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
X_15000_ net1206 vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__inv_2
XANTENNA__09766__B1 _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__B2 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ net1031 net1025 vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__nor2_1
XANTENNA__11995__B net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11573__A0 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12143_ net258 net2631 net511 vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_4__f_wb_clk_i clknet_3_2_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12117__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12074_ net242 net676 vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__and2_2
X_16951_ clknet_leaf_173_wb_clk_i _02620_ _01180_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10128__A1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ team_04_WB.MEM_SIZE_REG_REG\[24\] team_04_WB.MEM_SIZE_REG_REG\[23\] _06513_
+ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__or3_1
X_15902_ clknet_leaf_38_wb_clk_i _01579_ _00129_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__dfrtp_1
X_16882_ clknet_leaf_7_wb_clk_i _02551_ _01111_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\]
+ sky130_fd_sc_hd__dfrtp_1
X_15833_ clknet_leaf_90_wb_clk_i _01510_ _00060_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13078__A0 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15764_ net1284 vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__inv_2
XANTENNA__12825__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ net606 _07375_ net471 net315 net1816 vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a32o_1
X_14715_ net1126 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11927_ _03632_ _05955_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_157_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15695_ net1268 vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14646_ net1221 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ net652 net245 vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_99_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13250__A0 net87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _04357_ _04412_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14577_ net1260 vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11789_ net757 _05808_ net697 _03894_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12347__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ clknet_leaf_116_wb_clk_i _01985_ _00545_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[289\]
+ sky130_fd_sc_hd__dfrtp_1
X_13528_ team_04_WB.ADDR_START_VAL_REG\[22\] _02918_ vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_136_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17296_ net1352 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12066__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16247_ clknet_leaf_161_wb_clk_i _01916_ _00476_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[220\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13002__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] net1044 _02846_
+ net1081 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput115 net115 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__clkbuf_4
X_16178_ clknet_leaf_6_wb_clk_i _01847_ _00407_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput126 net126 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__clkbuf_4
XANTENNA__08655__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput137 net137 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15129_ net1251 vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__inv_2
Xoutput148 net148 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__12082__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput159 net159 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07951_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[18\] net1009
+ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_162_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07882_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] vssd1 vssd1
+ vccd1 vccd1 _03497_ sky130_fd_sc_hd__inv_2
XANTENNA__08732__A1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09621_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[99\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__mux2_1
XANTENNA__13608__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08719__B _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12816__A0 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[677\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[645\]
+ net951 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08503_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__inv_2
X_09483_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\]
+ net943 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11095__A2 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout255_A _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09862__A_N _04532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[824\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[792\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_1
XANTENNA__09330__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__A0 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ net642 _03974_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_1
XANTENNA__12044__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout422_A _07658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1164_A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08343__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13792__A1 _06932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08296_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout791_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout889_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_92 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_112_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1217_X net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout320 net321 vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_8
XANTENNA__13847__A2 _03235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 net332 vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_2
Xfanout342 net343 vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 _07484_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__clkbuf_8
Xfanout364 net365 vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout375 _07679_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__buf_2
XANTENNA__09071__S1 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 net387 vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_8
Xfanout397 _07670_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_4
X_09819_ _05426_ _05427_ _05428_ _05429_ net834 net746 vssd1 vssd1 vccd1 vccd1 _05430_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ _07528_ net327 net392 net1964 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a22o_1
XANTENNA__12807__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12761_ _07488_ net331 net398 net1784 vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__a22o_1
XANTENNA__12283__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14500_ net1285 vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__inv_2
X_11712_ _06709_ _06710_ _06861_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12692_ net2051 net405 net335 _07247_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a22o_1
X_15480_ net1205 vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13232__A0 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ team_04_WB.MEM_SIZE_REG_REG\[2\] _07090_ vssd1 vssd1 vccd1 vccd1 _07132_
+ sky130_fd_sc_hd__xnor2_1
X_14431_ net1291 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ clknet_leaf_85_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[4\]
+ _01379_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12586__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13783__B2 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14362_ net1262 vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11574_ net627 net589 net626 net580 net548 net542 vssd1 vssd1 vccd1 vccd1 _07063_
+ sky130_fd_sc_hd__mux4_2
Xinput17 DAT_I[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 DAT_I[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_1
X_16101_ clknet_leaf_169_wb_clk_i _01770_ _00330_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput39 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
X_13313_ net1083 team_04_WB.MEM_SIZE_REG_REG\[22\] team_04_WB.MEM_SIZE_REG_REG\[23\]
+ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__or3b_1
X_10525_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[25\]
+ _06088_ net1049 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14293_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\]
+ _03458_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__and3_1
X_17081_ clknet_leaf_45_wb_clk_i _00030_ _01310_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_165_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12338__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ net58 _06140_ _06146_ _06157_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__nand4_1
X_16032_ clknet_leaf_140_wb_clk_i _01701_ _00261_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ _06022_ _06031_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_131_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ _07611_ net375 net291 net1733 vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a22o_1
X_10387_ _05725_ _05742_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12126_ _06194_ _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__or2_1
X_16934_ clknet_leaf_21_wb_clk_i _02603_ _01163_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\]
+ sky130_fd_sc_hd__dfrtp_1
X_12057_ net822 _05279_ _04782_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__and3b_4
X_11008_ _06313_ _06493_ _06495_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09415__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A3 net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__B1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16865_ clknet_leaf_133_wb_clk_i _02534_ _01094_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_59 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15816_ clknet_leaf_89_wb_clk_i _01493_ _00043_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16796_ clknet_leaf_126_wb_clk_i _02465_ _01025_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15747_ net1275 vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _07627_ net473 net316 net1698 vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15678_ net1268 vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14629_ net1113 vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__inv_2
XANTENNA__12026__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_155_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13774__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12577__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08150_ net771 _03760_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08081_ _03686_ _03691_ net728 vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__mux2_1
X_17279_ net597 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
XANTENNA__08650__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11001__A2 _06489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__mux2_1
XANTENNA__09392__Y _05003_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07934_ net1051 _03543_ _03544_ _03535_ _03537_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__o221a_1
XANTENNA__09325__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12501__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A _07679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10698__C _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07921__X _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09535_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[389\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__mux2_1
XANTENNA__12265__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1281_A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__X _06932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\]
+ net889 vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08417_ _04010_ _04016_ _04027_ net716 vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a22o_2
X_09397_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[327\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12568__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08348_ _03955_ _03956_ _03957_ _03958_ net827 net744 vssd1 vssd1 vccd1 vccd1 _03959_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11776__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08279_ net772 _03883_ net765 vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__o21a_1
XFILLER_0_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10310_ net281 _05904_ net1056 vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11290_ _06279_ _06776_ _06778_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08619__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12434__B net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10241_ _05645_ net620 _05840_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a31o_1
XANTENNA__10235__A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05656_ _05780_ _05781_ net619 net281 vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1104 net1115 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__buf_4
Xfanout1115 net1158 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_2
XANTENNA__13480__A1_N net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1126 net1127 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__buf_4
X_14980_ net1189 vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__inv_2
Xfanout1137 net1138 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1148 net1150 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_4
Xfanout1159 net1166 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13931_ net132 net1072 net1041 _03297_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16650_ clknet_leaf_163_wb_clk_i _02319_ _00879_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\]
+ sky130_fd_sc_hd__dfrtp_1
X_13862_ _03226_ _03249_ net1809 net1066 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_87_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15601_ net1271 vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__inv_2
X_12813_ net251 net2629 net324 vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__mux2_1
X_16581_ clknet_leaf_185_wb_clk_i _02250_ _00810_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[554\]
+ sky130_fd_sc_hd__dfrtp_1
X_13793_ _07822_ _07823_ vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15532_ net1120 vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12744_ _07469_ net338 net401 net2057 vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09672__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15463_ net1141 vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__inv_2
XANTENNA__12008__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12675_ net253 net2389 net475 vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ net1408 _02812_ _01431_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14414_ net1277 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12559__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _05473_ _07107_ _07114_ net462 _07104_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o32a_2
XTAP_TAPCELL_ROW_133_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08662__X _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15394_ net1239 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08858__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ clknet_leaf_83_wb_clk_i team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[0\]
+ _01362_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14345_ net1190 vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__inv_2
X_11557_ net588 net547 _06574_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_40_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17064_ clknet_leaf_48_wb_clk_i _00011_ _01293_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10508_ _06077_ net1764 net1020 vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold609 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\] vssd1 vssd1
+ vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\]
+ _03447_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[20\] vssd1 vssd1
+ vccd1 vccd1 _03451_ sky130_fd_sc_hd__a31o_1
X_11488_ _06383_ _06427_ _06381_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17196__Q team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_562 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09188__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16015_ clknet_leaf_53_wb_clk_i _01691_ _00244_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13227_ net74 team_04_WB.MEM_SIZE_REG_REG\[14\] net983 vssd1 vssd1 vccd1 vccd1 _01676_
+ sky130_fd_sc_hd__mux2_1
X_10439_ _06009_ _06014_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12731__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _07594_ net376 net292 net2016 vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__a22o_1
XANTENNA__10742__A1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13456__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ net1996 net354 _07509_ net450 vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__a22o_1
X_13089_ net699 _05279_ _06181_ _07666_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__or4_4
X_16917_ clknet_leaf_34_wb_clk_i _02586_ _01146_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\]
+ sky130_fd_sc_hd__dfrtp_1
X_16848_ clknet_leaf_191_wb_clk_i _02517_ _01077_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08984__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12247__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16779_ clknet_leaf_15_wb_clk_i _02448_ _01008_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[752\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12359__X _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13191__A _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[168\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[136\]
+ net957 vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__mux2_1
XANTENNA__09112__B2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13995__A1 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _04858_ _04859_ _04860_ _04861_ net824 net741 vssd1 vssd1 vccd1 vccd1 _04862_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_168_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08202_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[509\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09182_ net722 _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_170_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08133_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[542\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_170_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout218_A _07277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net973 _03673_ vssd1 vssd1 vccd1
+ vccd1 _03675_ sky130_fd_sc_hd__o21ai_4
XANTENNA__08224__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12254__B net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14750__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09274__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1127_A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12722__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10733__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A _05139_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12270__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[623\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[591\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__mux2_1
X_07917_ _03527_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout754_A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08897_ net722 _04507_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__or2_1
XANTENNA__10497__B1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15581__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08894__S net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_162_Right_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09518_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[932\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[900\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790_ net466 _06278_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nor2_2
XFILLER_0_151_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[326\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12460_ net519 net600 _07461_ net428 net1959 vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a32o_1
XANTENNA__11749__A0 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11411_ net755 _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12391_ _07445_ net2373 net498 vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14130_ team_04_WB.MEM_SIZE_REG_REG\[29\] _07703_ _07706_ team_04_WB.ADDR_START_VAL_REG\[29\]
+ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__a22o_1
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11342_ _06788_ _06796_ net562 vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__mux2_1
XANTENNA__12961__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11273_ team_04_WB.MEM_SIZE_REG_REG\[17\] _06509_ vssd1 vssd1 vccd1 vccd1 _06762_
+ sky130_fd_sc_hd__xnor2_1
X_14061_ net24 net1063 _03352_ team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1
+ vccd1 vccd1 _01525_ sky130_fd_sc_hd__a22o_1
XANTENNA__14660__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08917__A1 net661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input50_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ net620 _05827_ net277 vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_37_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12713__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ net602 _07472_ net469 net310 net1981 vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_37_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08393__A2 _04002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _05680_ _05681_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09017__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _04559_ vssd1
+ vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__or2_1
XANTENNA__11508__B _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ net1232 vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold6 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\] vssd1 vssd1 vccd1
+ vccd1 net1443 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13674__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output137_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ clknet_leaf_142_wb_clk_i _02371_ _00931_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ _02991_ _03278_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_8 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14894_ net1195 vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_50_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16633_ clknet_leaf_177_wb_clk_i _02302_ _00862_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\]
+ sky130_fd_sc_hd__dfrtp_1
X_13845_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[31\] net1044 _03235_
+ net1081 net1002 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__o221a_1
XANTENNA__12229__B2 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13977__B2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16564_ clknet_leaf_3_wb_clk_i _02233_ _00793_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13776_ net709 _03160_ _03163_ net998 _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10988_ _06352_ _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12339__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15515_ net1138 vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _07452_ net340 net402 net1957 vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__a22o_1
X_16495_ clknet_leaf_186_wb_clk_i _02164_ _00724_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10660__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ net1223 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__inv_2
X_12658_ net218 net2625 net476 vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11609_ _07013_ _07097_ net563 vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15377_ net1276 vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12589_ _07558_ net481 net412 net1901 vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XANTENNA__12355__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__B2 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17116_ clknet_leaf_105_wb_clk_i _02751_ _01345_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14328_ _03519_ _03484_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12074__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold406 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[418\] vssd1 vssd1
+ vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\] vssd1 vssd1
+ vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold428 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[121\] vssd1 vssd1
+ vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17047_ clknet_leaf_173_wb_clk_i _02716_ _01276_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_78_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold439 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\] vssd1 vssd1
+ vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14259_ net1807 _03438_ _03440_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08979__S net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12704__A2 net405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout908 net910 vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_4
Xfanout919 net920 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_74_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _04427_ _04428_ _04429_ _04430_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04431_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09581__A1 _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_146_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\] vssd1 vssd1
+ vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\] vssd1 vssd1
+ vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
Xhold1128 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[895\] vssd1 vssd1
+ vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1139 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[398\] vssd1 vssd1
+ vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_124_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07912__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09603__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08219__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_424 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09303_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[713\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_172_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12640__A1 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14745__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_124_wb_clk_i_A clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_91_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ _04841_ _04842_ _04843_ _04844_ net824 net741 vssd1 vssd1 vccd1 vccd1 _04845_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[523\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_A _07591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1244_A net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08116_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[30\] team_04_WB.instance_to_wrap.CPU_DAT_O\[30\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__mux2_2
XANTENNA__10403__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[141\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13795__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] net1079 net1028 net1024 vssd1
+ vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12156__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[579\] vssd1 vssd1
+ vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08889__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14480__A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold951 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[863\] vssd1 vssd1
+ vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\] vssd1 vssd1
+ vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[421\] vssd1 vssd1
+ vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[67\] vssd1 vssd1
+ vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[773\] vssd1 vssd1
+ vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout871_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout969_A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ net625 _05282_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_32_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[79\]
+ net897 vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__mux2_1
XANTENNA__12459__B2 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09324__A1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ net2354 net528 net451 _07421_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_163_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_174_Left_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ net588 _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nor2_1
X_11891_ net655 net256 vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__and2_1
X_13630_ net993 _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13959__A1 _03918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10842_ _03946_ _06329_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _05904_ net1100
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10773_ net644 net550 _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15300_ net1169 vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__inv_2
X_12512_ _07509_ net487 net426 net1838 vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16280_ clknet_leaf_156_wb_clk_i _01949_ _00509_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[253\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input98_A wbs_dat_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ net997 _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13187__A2 net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15231_ net1250 vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__inv_2
XANTENNA__11350__Y _06839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10394__S net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12443_ net2512 net430 _07642_ net523 vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08063__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15162_ net1137 vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__inv_2
X_12374_ net244 net2419 net498 vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ team_04_WB.MEM_SIZE_REG_REG\[12\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[12\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__o221a_4
XFILLER_0_120_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11325_ _06279_ _06808_ _06813_ _04248_ _06812_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__a221o_1
X_15093_ net1211 vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__inv_2
XANTENNA__12147__A0 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08799__S net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14044_ net12 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1 vssd1
+ vccd1 vccd1 _01542_ sky130_fd_sc_hd__a22o_1
X_11256_ _06547_ _06587_ net553 vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
XANTENNA__09012__B1 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13895__B1 _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09915__C net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ net619 _05810_ _05812_ net280 vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a211o_1
XANTENNA__08997__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11187_ _06272_ _06674_ _06675_ net585 vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10138_ _05715_ _05748_ _05716_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__o21a_1
X_15995_ clknet_leaf_70_wb_clk_i _01671_ _00224_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13647__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11806__X _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13111__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[23\] _04113_ vssd1
+ vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__or2_1
X_14946_ net1265 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11122__A1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14877_ net1155 vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16616_ clknet_leaf_113_wb_clk_i _02285_ _00845_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\]
+ sky130_fd_sc_hd__dfrtp_1
X_13828_ team_04_WB.ADDR_START_VAL_REG\[24\] _03218_ vssd1 vssd1 vccd1 vccd1 _03219_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_148_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16547_ clknet_leaf_124_wb_clk_i _02216_ _00776_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[520\]
+ sky130_fd_sc_hd__dfrtp_1
X_13759_ _07827_ _07829_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11830__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16478_ clknet_leaf_115_wb_clk_i _02147_ _00707_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_54 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15429_ net1109 vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__inv_2
XANTENNA__13178__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12386__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11189__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold203 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[11\] vssd1
+ vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold214 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\] vssd1 vssd1
+ vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_76_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 net134 vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A0 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\] vssd1 vssd1
+ vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold247 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\] vssd1 vssd1
+ vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\] vssd1 vssd1
+ vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\] team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[12\]
+ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__and3_1
XANTENNA__09394__A _03724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold269 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\] vssd1 vssd1
+ vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09003__B1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout705 _03632_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11429__A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout716 _03674_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_165_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__C1 net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ net698 _05451_ _03621_ net905 vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__and4b_2
Xfanout727 net728 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__clkbuf_8
Xfanout738 net739 vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_165_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 net750 vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__buf_2
X_08803_ net591 _04412_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__xnor2_1
X_09783_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\]
+ net961 vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__mux2_1
XANTENNA__10052__B _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13644__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\]
+ net868 vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
XANTENNA__09333__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1194_A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08596_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\]
+ net908 vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout717_A _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13169__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09217_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12377__A0 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__C net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[11\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14118__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14118__B2 team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__B2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
XANTENNA__12129__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ _03865_ net364 net360 _03863_ _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__o221a_1
Xclkbuf_4_3__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_12090_ net259 net677 vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_9_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08412__S net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\] vssd1 vssd1
+ vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold781 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[590\] vssd1 vssd1
+ vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold792 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\] vssd1 vssd1
+ vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net566 _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14800_ net1165 vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__inv_2
XANTENNA__11626__X _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15780_ net1259 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__inv_2
X_12992_ _07643_ net473 net312 net2010 vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09243__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input13_A DAT_I[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ net1161 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__inv_2
X_11943_ _07398_ _07406_ _07405_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__a21oi_1
X_14662_ net1106 vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__inv_2
X_11874_ _06920_ _06931_ net689 vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16401_ clknet_leaf_179_wb_clk_i _02070_ _00630_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[374\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13613_ net1001 _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10825_ _03721_ _06312_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__and2_1
X_14593_ net1182 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11802__A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16332_ clknet_leaf_120_wb_clk_i _02001_ _00561_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[305\]
+ sky130_fd_sc_hd__dfrtp_1
X_13544_ _07830_ _07833_ _07835_ _07839_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10756_ _06242_ _06244_ net530 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16263_ clknet_leaf_22_wb_clk_i _01932_ _00492_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\]
+ sky130_fd_sc_hd__dfrtp_1
X_13475_ _07859_ _07862_ _07865_ _07869_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__or4_1
X_10687_ net1701 net711 _06180_ net2326 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09459__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15214_ net1204 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12426_ net654 net608 net233 vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__and3_1
XANTENNA__12907__A2 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16194_ clknet_leaf_143_wb_clk_i _01863_ _00423_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11948__S _07234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15145_ net1133 vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__inv_2
X_12357_ _07443_ _07444_ net671 vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__and3_2
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _06581_ _06584_ net539 vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__mux2_1
X_15076_ net1171 vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__inv_2
X_12288_ net228 net674 vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__and2_1
X_14027_ net2004 net1068 net1039 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__a21o_1
XANTENNA__11879__C1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11239_ net286 _06723_ _06725_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_143_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09942__A _03892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15978_ clknet_leaf_52_wb_clk_i _01654_ _00207_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_160_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14929_ net1267 vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08450_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[440\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15800__19 clknet_leaf_61_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__inv_2
X_08381_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[985\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11803__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12071__A2 net353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09002_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[334\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_115_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13639__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__S1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_158_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_158_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_167_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10385__A2 net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09328__S net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08232__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__B net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ _05502_ _05504_ _05506_ _04088_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 _07591_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout513 net514 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__buf_6
Xfanout524 net525 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout535 net536 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_2
Xfanout546 _05377_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
X_09835_ _03621_ _05441_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__nand3_2
Xfanout557 net558 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
XANTENNA_input5_A DAT_I[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout568 _05251_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__buf_2
XANTENNA__11885__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 _05219_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_2
XANTENNA_fanout667_A _03633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09766_ net664 _05375_ _05340_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09063__S net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ net765 _04321_ _04327_ _04315_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__a31oi_4
XANTENNA__08189__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__B _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ net667 _05283_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout455_X net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08648_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[53\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[21\]
+ net907 vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13821__B net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08579_ _04186_ _04187_ _04188_ _04189_ net825 net742 vssd1 vssd1 vccd1 vccd1 _04190_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12598__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09689__S1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ net44 net43 net46 net45 vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__or4b_1
XFILLER_0_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11590_ _06414_ _07078_ net462 vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__B1 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ _06099_ net2024 net1022 vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13260_ net76 team_04_WB.ADDR_START_VAL_REG\[16\] net975 vssd1 vssd1 vccd1 vccd1
+ _01646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13011__A1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ _03531_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09215__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ net233 net649 vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13191_ _06174_ net1001 vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11573__A1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09238__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12142_ net259 net2630 net512 vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
XANTENNA__08142__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12073_ net2219 net352 _07491_ net436 vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
X_16950_ clknet_leaf_12_wb_clk_i _02619_ _01179_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\]
+ sky130_fd_sc_hd__dfrtp_1
X_11024_ team_04_WB.MEM_SIZE_REG_REG\[22\] _06512_ vssd1 vssd1 vccd1 vccd1 _06513_
+ sky130_fd_sc_hd__or2_1
X_15901_ clknet_leaf_38_wb_clk_i _01578_ _00128_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__dfrtp_1
XANTENNA__09762__A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16881_ clknet_leaf_176_wb_clk_i _02550_ _01110_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\]
+ sky130_fd_sc_hd__dfrtp_1
X_15832_ clknet_leaf_91_wb_clk_i _01509_ _00059_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10701__A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15763_ net1283 vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
X_12975_ net610 _07369_ net474 net317 net1680 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a32o_1
XANTENNA__10420__B net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14714_ net1146 vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__inv_2
X_11926_ team_04_WB.instance_to_wrap.CPU_DAT_O\[8\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07392_ sky130_fd_sc_hd__a21o_1
XANTENNA__14027__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15694_ net1268 vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14645_ net1207 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__inv_2
X_11857_ net689 _06757_ _07332_ net613 vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__o211a_2
XFILLER_0_170_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14319__S net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12589__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ _04474_ _04528_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__and2_1
X_14576_ net1260 vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08317__S net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11788_ team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07273_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12347__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16315_ clknet_leaf_103_wb_clk_i _01984_ _00544_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[288\]
+ sky130_fd_sc_hd__dfrtp_1
X_13527_ net709 _02911_ _02914_ net996 _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_136_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17295_ net1351 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_166_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10739_ _06227_ net646 _06226_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_136_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16246_ clknet_leaf_15_wb_clk_i _01915_ _00475_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13458_ _07691_ _02848_ _02847_ net1002 vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a211o_1
XANTENNA__13002__A1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ net2153 net432 _07632_ net520 vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
XANTENNA__10582__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16177_ clknet_leaf_172_wb_clk_i _01846_ _00406_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__clkbuf_4
X_13389_ _07769_ _07813_ _07814_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput116 net116 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput127 net127 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12761__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15128_ net1203 vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__inv_2
Xoutput138 net138 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput149 net149 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12082__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07950_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[319\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__mux2_1
X_15059_ net1244 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_162_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12513__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[26\] vssd1 vssd1
+ vccd1 vccd1 _03496_ sky130_fd_sc_hd__inv_2
XANTENNA__11867__A2 net529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__mux2_1
X_09551_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[741\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\]
+ net951 vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08502_ net751 net729 _03725_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__a21o_2
X_09482_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\]
+ net946 vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08433_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[856\]
+ net916 vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout248_A _07307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12044__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08227__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08343__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13792__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08295_ net729 _03905_ net713 vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1157_A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09058__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__Y _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 _07678_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_4
XANTENNA__12504__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout321 _07675_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_4
Xfanout332 _07667_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_2
Xfanout343 net351 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout354 net355 vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08184__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _06249_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
Xfanout376 net377 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__clkbuf_4
X_09818_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[897\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__mux2_1
Xfanout387 _07674_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10521__A team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout398 _07670_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08198__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09359__S0 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09749_ _05356_ _05357_ _05358_ _05359_ net837 net739 vssd1 vssd1 vccd1 vccd1 _05360_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10818__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ _07487_ net340 net398 net1687 vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__a22o_1
XANTENNA__12283__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13480__B2 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_6_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09521__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11711_ _06655_ _06656_ _07169_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12691_ _06189_ net614 _06196_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__and3b_4
XFILLER_0_51_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12448__A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14430_ net1277 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__inv_2
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11642_ _07119_ _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08137__S net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12167__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ net1262 vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ net626 net580 net548 vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 DAT_I[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ clknet_leaf_168_wb_clk_i _01769_ _00329_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input80_A wbs_dat_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ net1083 team_04_WB.MEM_SIZE_REG_REG\[22\] vssd1 vssd1 vccd1 vccd1 _07738_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12991__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ clknet_leaf_45_wb_clk_i _00028_ _01309_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput29 DAT_I[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] net1096 net1051 vssd1 vssd1 vccd1
+ vccd1 _06088_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_94_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14292_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[24\]
+ _03457_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[26\] vssd1 vssd1
+ vccd1 vccd1 _03461_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16031_ clknet_leaf_155_wb_clk_i _01700_ _00260_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_13243_ net58 _06146_ _06152_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__nand3_1
XFILLER_0_161_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10455_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _06032_
+ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__nor2_1
XFILLER_0_161_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12183__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10349__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12743__B1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _07610_ net377 net292 net1607 vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a22o_1
X_10386_ _05603_ _05604_ _05618_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _05221_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09763__Y _05374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ net2601 net518 _07481_ net460 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a22o_1
X_16933_ clknet_leaf_170_wb_clk_i _02602_ _01162_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_9__f_wb_clk_i_A clknet_3_4_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13218__S net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _06313_ _06493_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__or3_1
X_16864_ clknet_leaf_136_wb_clk_i _02533_ _01093_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\]
+ sky130_fd_sc_hd__dfrtp_1
X_15815_ clknet_leaf_77_wb_clk_i _01492_ _00042_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_16795_ clknet_leaf_96_wb_clk_i _02464_ _01024_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15746_ net1294 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _07626_ net473 net316 net1818 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11909_ net760 _05934_ net695 _07377_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_138_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15677_ net1281 vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__inv_2
XFILLER_0_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12889_ _05221_ _07590_ _07663_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__or3_4
XFILLER_0_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14628_ net1167 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__inv_2
XANTENNA__13223__A1 team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12026__A2 net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14559_ net1182 vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__inv_2
XANTENNA__12792__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14573__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _03687_ _03688_ _03689_ _03690_ net827 net743 vssd1 vssd1 vccd1 vccd1 _03691_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12982__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17278_ team_04_WB.instance_to_wrap.final_design.pixel_data vssd1 vssd1 vccd1 vccd1
+ net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08650__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ clknet_leaf_4_wb_clk_i _01898_ _00458_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12734__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08982_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[174\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[142\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_143_Right_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07933_ net1051 _03543_ _03544_ _03535_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__o22ai_1
XANTENNA__09589__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[675\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10060__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_155_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09534_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[485\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[453\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09666__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09341__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _05072_ _05073_ _05074_ _05075_ net835 net745 vssd1 vssd1 vccd1 vccd1 _05076_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09761__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12268__A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1274_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08416_ _04021_ _04026_ net720 vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__mux2_1
X_09396_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\]
+ net878 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11225__A0 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09513__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_173_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_173_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout320_X net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08347_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[442\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12973__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_102_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ net778 _03888_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout999_A _07686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12725__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ net620 _05841_ net277 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__A1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _05664_ _05774_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1107 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_4
XANTENNA__09516__S net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1116 net1118 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1127 net1158 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1138 net1157 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_2
Xfanout1149 net1150 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_4
XANTENNA__13150__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _03097_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_35_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13861_ _02875_ _03225_ net1039 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_87_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14658__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15600_ net1163 vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12812_ _07385_ net2543 net322 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__mux2_1
X_16580_ clknet_leaf_171_wb_clk_i _02249_ _00809_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\]
+ sky130_fd_sc_hd__dfrtp_1
X_13792_ _06932_ net272 net710 vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a21o_1
X_15531_ net1159 vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__inv_2
XFILLER_0_167_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12743_ _07468_ net346 net403 net1963 vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ net1104 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12008__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12674_ net254 net2467 net475 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17201_ clknet_leaf_78_wb_clk_i team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[1\]
+ _01430_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ net1274 vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _06776_ _06948_ _07110_ _07111_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__a221o_1
XANTENNA__11216__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12__f_wb_clk_i_X clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15393_ net1129 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11767__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ clknet_leaf_66_wb_clk_i _02767_ _01361_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12964__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14344_ net1190 vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__inv_2
XANTENNA_input83_X net83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11556_ net626 net547 net541 _06579_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__a211o_1
XANTENNA__08632__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17063_ clknet_leaf_49_wb_clk_i _00010_ _01292_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10507_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[31\]
+ _06076_ net1047 vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14275_ net1945 _03448_ _03450_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_150_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11487_ _06973_ _06974_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16014_ clknet_leaf_47_wb_clk_i _01690_ _00243_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12716__B1 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__B2 net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ net75 team_04_WB.MEM_SIZE_REG_REG\[15\] net982 vssd1 vssd1 vccd1 vccd1 _01677_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10438_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[3\] _06016_
+ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11956__S net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12192__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ _07593_ net371 net290 net1836 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__a22o_1
XANTENNA__11419__A1_N net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10369_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] net1057 vssd1
+ vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12108_ _07402_ net678 vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__and2_1
XANTENNA__13456__B _02846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13088_ _07445_ net2494 net305 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__mux2_1
XANTENNA__13141__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16916_ clknet_leaf_2_wb_clk_i _02585_ _01145_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\]
+ sky130_fd_sc_hd__dfrtp_1
X_12039_ net249 net684 vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__and2_1
XANTENNA__12495__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16847_ clknet_leaf_189_wb_clk_i _02516_ _01076_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14568__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12247__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778_ clknet_leaf_166_wb_clk_i _02447_ _01007_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13191__B net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15729_ net1295 vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13995__A2 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12088__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_114_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09250_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[682\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[650\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08201_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\]
+ net943 vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ _04788_ _04789_ _04790_ _04791_ net828 net735 vssd1 vssd1 vccd1 vccd1 _04792_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12955__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08132_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[638\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[606\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_78_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_170_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10607__Y _06145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08063_ team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] net973 _03673_ vssd1 vssd1 vccd1
+ vccd1 _03674_ sky130_fd_sc_hd__o21a_4
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12970__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12707__B1 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10055__B _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1022_A _06073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08240__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _04572_ _04573_ _04574_ _04575_ net831 net747 vssd1 vssd1 vccd1 vccd1 _04576_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12270__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout482_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_87_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08896_ _04503_ _04504_ _04505_ _04506_ net829 net744 vssd1 vssd1 vccd1 vccd1 _04507_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12486__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_153_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10497__B2 team_04_WB.instance_to_wrap.final_design.VGA_adr\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8__f_wb_clk_i_X clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09517_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11614__B _07102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout914_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09448_ net667 _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_96_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ net780 _04989_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__or2_1
XANTENNA__12946__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ net462 _06883_ _06898_ _05473_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__o22a_1
X_12390_ _07438_ net2572 net498 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11341_ net573 _06826_ _06828_ _06829_ net586 vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14060_ net27 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1
+ vccd1 vccd1 _01526_ sky130_fd_sc_hd__a22o_1
X_11272_ _06758_ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08378__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12174__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ net601 _07471_ net468 net310 net1710 vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a32o_1
X_10223_ _05679_ _05767_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08917__A2 _04526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_192_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10185__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11921__A1 _03631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__B2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10154_ _05683_ _05764_ _05682_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_89_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13123__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ net1238 vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__inv_2
X_10085_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] _04502_ vssd1
+ vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__xnor2_1
Xhold7 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[30\] vssd1 vssd1 vccd1
+ vccd1 net1444 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12477__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__B2 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ clknet_leaf_131_wb_clk_i _02370_ _00930_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13913_ net1859 net1071 net1040 _03285_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__a22o_1
XANTENNA__11685__B1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14893_ net1152 vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13844_ _03233_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__xnor2_2
X_16632_ clknet_leaf_149_wb_clk_i _02301_ _00861_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[605\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13426__A1 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12229__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13775_ net1002 _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__or2_1
XANTENNA__13977__A2 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16563_ clknet_leaf_183_wb_clk_i _02232_ _00792_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ net638 _06351_ _06348_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__o21a_1
XFILLER_0_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12726_ _07451_ net340 net402 net2002 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__a22o_1
X_15514_ net1151 vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16494_ clknet_leaf_27_wb_clk_i _02163_ _00723_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[467\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ net1209 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10660__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_12657_ net220 net2312 net475 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__mux2_1
XANTENNA__13231__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12937__A0 _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ _07062_ _07096_ net542 vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ net1162 vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12588_ _07557_ net483 net413 net2150 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12401__A2 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12355__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14327_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[3\] _03483_
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] _03520_ vssd1
+ vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17115_ clknet_leaf_91_wb_clk_i _02750_ _01344_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11539_ net628 net627 net589 net626 net547 net541 vssd1 vssd1 vccd1 vccd1 _07028_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold407 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[97\] vssd1 vssd1
+ vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold418 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[380\] vssd1 vssd1
+ vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ clknet_leaf_11_wb_clk_i _02715_ _01275_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
X_14258_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] _03438_
+ net820 vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__o21ai_1
Xhold429 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[629\] vssd1 vssd1
+ vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_78_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13209_ net61 _06140_ _06145_ _06158_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nand4_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09030__A1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14189_ _03530_ _03374_ _03380_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.v_out
+ sky130_fd_sc_hd__or3b_1
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__B net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[306\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[274\]
+ net933 vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__mux2_1
Xhold1107 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\] vssd1 vssd1
+ vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08216__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1118 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[791\] vssd1 vssd1
+ vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08995__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1129 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[134\] vssd1 vssd1
+ vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12468__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ _04288_ _04289_ _04290_ _04291_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04292_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11715__A _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_84 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__A1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[553\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_172_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12640__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[394\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10651__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout230_A _07426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12928__A0 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout328_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09164_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__mux2_1
XANTENNA__08235__S net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _03639_ _03641_ _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__a21o_4
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09095_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[237\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[205\]
+ net963 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1237_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1126 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_2__f_wb_clk_i clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
X_08046_ net1008 net1007 vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold930 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\] vssd1 vssd1
+ vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[484\] vssd1 vssd1
+ vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold952 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[522\] vssd1 vssd1
+ vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[971\] vssd1 vssd1
+ vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold974 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\] vssd1 vssd1
+ vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[867\] vssd1 vssd1
+ vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\] vssd1 vssd1
+ vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _05606_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13105__B1 net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _03554_ net703 _04330_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a21o_1
XANTENNA__12459__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15806__25 clknet_leaf_55_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout652_X net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__mux2_1
X_10910_ net583 _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13408__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ net695 _07150_ _07361_ net615 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a211oi_2
XANTENNA__14001__A _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13959__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ net642 _06329_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout917_X net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13560_ net1093 _02950_ net1044 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__o2bb2a_1
X_10772_ net643 net550 vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_1
XANTENNA__08835__A1 _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12631__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12511_ _07508_ net492 net427 net1998 vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ net994 _02878_ _02881_ _07691_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a22o_1
XANTENNA__12456__A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12919__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15230_ net1214 vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12442_ net607 net213 net682 vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12175__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13592__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ net1251 vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__inv_2
X_12373_ net245 net2610 net496 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14671__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ team_04_WB.MEM_SIZE_REG_REG\[11\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[11\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__o221a_4
X_11324_ _04247_ _06248_ net362 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a21o_1
X_15092_ net1214 vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14043_ net14 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1
+ vccd1 vccd1 _01543_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_56_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09012__A1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ net582 _06743_ net288 vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__o21a_1
XANTENNA__12191__A _07349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12698__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ net619 _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_128_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08997__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _06555_ _06588_ net567 vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10137_ _05745_ _05747_ _05717_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__a21oi_1
X_15994_ clknet_leaf_71_wb_clk_i _01670_ _00223_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09704__S net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ _05677_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14945_ net1188 vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__inv_2
XANTENNA__11535__A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12130__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15007__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10330__B1 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14876_ net1128 vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__inv_2
XANTENNA__12870__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16615_ clknet_leaf_165_wb_clk_i _02284_ _00844_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\]
+ sky130_fd_sc_hd__dfrtp_1
X_13827_ net709 _03212_ _03214_ net996 _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_723 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17299__1355 vssd1 vssd1 vccd1 vccd1 _17299__1355/HI net1355 sky130_fd_sc_hd__conb_1
XFILLER_0_159_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14846__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ net753 _06729_ net272 net709 vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_98 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16546_ clknet_leaf_147_wb_clk_i _02215_ _00775_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12622__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12709_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\] net407 net347
+ _07363_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10585__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11830__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ team_04_WB.ADDR_START_VAL_REG\[1\] _03073_ vssd1 vssd1 vccd1 vccd1 _03080_
+ sky130_fd_sc_hd__xor2_1
X_16477_ clknet_leaf_127_wb_clk_i _02146_ _00706_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15428_ net1171 vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15359_ net1249 vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__inv_2
XANTENNA__12653__X _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold204 net117 vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14127__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold215 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\] vssd1 vssd1
+ vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold226 net126 vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[317\] vssd1 vssd1
+ vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
X_09920_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[11\] _05530_ vssd1
+ vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__and2_1
Xhold248 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[255\] vssd1 vssd1
+ vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 net106 vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09394__B _03893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17029_ clknet_leaf_185_wb_clk_i _02698_ _01258_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08437__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout706 net707 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__clkbuf_4
Xfanout717 _03674_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
X_09851_ net698 _05451_ _03621_ net905 vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__nand4b_2
XFILLER_0_1_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11429__B _06915_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 net732 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_165_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _03649_ vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
X_08802_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__inv_2
X_09782_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\]
+ net961 vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09614__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07923__A _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12310__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08664_ _04274_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__inv_2
XANTENNA__12861__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08595_ net770 _04199_ net761 vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout445_A net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14063__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13810__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08754__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12613__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12276__A net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[842\]
+ net922 vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_699 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09147_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[107\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14118__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[844\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08029_ _03615_ _03622_ _03635_ _03637_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__or4_4
XFILLER_0_13_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10524__A team_04_WB.instance_to_wrap.CPU_DAT_O\[25\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold760 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[821\] vssd1 vssd1
+ vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\] vssd1 vssd1
+ vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12442__C net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[953\] vssd1 vssd1
+ vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ net558 net536 _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__nand4_1
Xhold793 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\] vssd1 vssd1
+ vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12991_ _07642_ net473 net312 net2212 vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11942_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[6\] team_04_WB.instance_to_wrap.CPU_DAT_O\[6\]
+ _07234_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14730_ net1106 vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10312__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08600__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12852__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14661_ net1113 vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__inv_2
X_11873_ net687 _07346_ _07343_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14054__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13612_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[7\] net1045 _02996_
+ net1098 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a2bb2o_1
X_16400_ clknet_leaf_192_wb_clk_i _02069_ _00629_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10824_ _03721_ _06312_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__nor2_1
X_14592_ net1185 vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08664__A _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12604__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09112__X _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13543_ _06816_ net272 net709 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16331_ clknet_leaf_23_wb_clk_i _02000_ _00560_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ net595 net549 _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11090__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ clknet_leaf_19_wb_clk_i _01931_ _00491_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\]
+ sky130_fd_sc_hd__dfrtp_1
X_13474_ _07166_ net273 _07697_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__o21ai_1
X_10686_ net2326 net711 _06180_ net2591 vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output197_A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15213_ net1199 vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12425_ net523 net607 _07403_ net434 net1634 vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_97_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16193_ clknet_leaf_141_wb_clk_i _01862_ _00422_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[166\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14109__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ net1125 vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__inv_2
X_12356_ net2275 net501 _07622_ net455 vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__a22o_1
XANTENNA__08603__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11307_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__inv_2
X_15075_ net1165 vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12287_ net2539 net505 _07586_ net455 vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
XANTENNA__13868__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ net1463 net1072 _03307_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__a21bo_1
X_11238_ _04359_ net363 net360 _04358_ _06726_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_71_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11879__B1 _06184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12540__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11817__X _07298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09942__B _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _06476_ _06657_ _06345_ _06352_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15977_ clknet_leaf_43_wb_clk_i _01653_ _00206_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13096__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14928_ net1173 vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12843__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15797__16 clknet_leaf_60_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__inv_2
XANTENNA__12795__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14859_ net1167 vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__inv_2
XANTENNA__14045__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[825\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[793\]
+ net906 vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11803__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16529_ clknet_leaf_179_wb_clk_i _02198_ _00758_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12096__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09472__B2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ net703 _04611_ _04386_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15200__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08432__C1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09903_ _03920_ _03977_ _05513_ _05512_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__a31o_1
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout514 _07519_ vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_4
XFILLER_0_10_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout525 _06197_ vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_4
XANTENNA_fanout395_A _07672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout536 net538 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
X_09834_ _04669_ _04725_ _04611_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a21o_4
Xclkbuf_leaf_127_wb_clk_i clknet_4_11__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout547 net548 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
XANTENNA__14103__X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 _05309_ vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_2
Xfanout569 _05251_ vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_4
X_09765_ net664 _05375_ _05340_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08716_ net778 _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__or2_1
X_09696_ net719 _05306_ _05295_ _05294_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12834__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A3 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08647_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[117\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[85\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14036__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout827_A net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[694\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11270__A1 team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[20\]
+ _06098_ net1049 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _06037_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__nand2_1
XANTENNA__09215__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_157_Right_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08649__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__C1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ net2448 net509 _07546_ net453 vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13190_ _06175_ net1001 vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_2
XANTENNA__08423__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09766__A2 _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ net244 net2369 net514 vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17298__1354 vssd1 vssd1 vccd1 vccd1 _17298__1354/HI net1354 sky130_fd_sc_hd__conb_1
XFILLER_0_124_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ net226 net676 vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__and2_1
Xhold590 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\] vssd1 vssd1
+ vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__A1 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13565__A team_04_WB.ADDR_START_VAL_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ team_04_WB.MEM_SIZE_REG_REG\[21\] team_04_WB.MEM_SIZE_REG_REG\[20\] _06511_
+ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__or3_1
X_15900_ clknet_leaf_120_wb_clk_i _01577_ _00127_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__dfrtp_1
X_16880_ clknet_leaf_192_wb_clk_i _02549_ _01109_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15831_ clknet_leaf_93_wb_clk_i _01508_ _00058_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_32_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15780__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11085__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15762_ net1269 vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__inv_2
X_12974_ net611 _07363_ net474 net317 net1591 vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__a32o_1
XANTENNA__12825__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14713_ net1238 vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__inv_2
X_11925_ net1983 net526 net442 _07391_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a22o_1
XANTENNA__14396__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15693_ net1267 vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ net686 _07331_ _07330_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__a21o_1
X_14644_ net1208 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_99_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ net658 _06291_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_99_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ net1260 vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__inv_2
X_11787_ net2005 net526 net441 _07272_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08888__S0 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16314_ clknet_leaf_44_wb_clk_i _01983_ _00543_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[287\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13526_ net996 _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nand2_1
X_10738_ net569 _05446_ net467 _05469_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__or4_2
X_17294_ net1350 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_136_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13457_ _03493_ _05784_ net1100 vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__mux2_1
X_16245_ clknet_leaf_32_wb_clk_i _01914_ _00474_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\]
+ sky130_fd_sc_hd__dfrtp_1
X_10669_ net1578 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[12\] vssd1
+ vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09429__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ net652 net602 net247 vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__and3_1
XFILLER_0_141_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13388_ _07769_ _07812_ _07806_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__a21o_1
X_16176_ clknet_leaf_3_wb_clk_i _01845_ _00405_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput117 net117 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__clkbuf_4
XANTENNA__12761__A1 _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput128 net128 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__clkbuf_4
X_15127_ net1230 vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__inv_2
X_12339_ net251 net668 vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__and2_2
Xoutput139 net139 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09953__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15058_ net1244 vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09065__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14009_ net1438 net1069 _03340_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a21o_1
X_07880_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] vssd1 vssd1
+ vccd1 vccd1 _03495_ sky130_fd_sc_hd__inv_2
XANTENNA__14070__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_50_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09164__S net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07940__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09550_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[549\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08501_ net766 _04111_ _04100_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_108_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09481_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[228\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\]
+ net945 vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08432_ net779 _04042_ _04037_ net761 vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08363_ net663 _03973_ _03949_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10339__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ _03901_ _03902_ _03903_ _03904_ net828 net735 vssd1 vssd1 vccd1 vccd1 _03905_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_A _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A _07661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09339__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout311 _07678_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout398_X net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 _07671_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_6
Xfanout333 net337 vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__clkbuf_4
Xfanout344 net345 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_4
Xfanout355 _07484_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_4
XANTENNA__08184__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09074__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__mux2_1
Xfanout377 net381 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_4
Xfanout388 _07673_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_6
XANTENNA__10521__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 _07670_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09359__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\]
+ net903 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11904__Y _07374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[290\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[258\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__mux2_1
XANTENNA__09684__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11192__X _06681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11710_ _06523_ _06592_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_95_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15105__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12690_ net610 _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__nor2_4
XANTENNA__08418__S net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11641_ net755 _07129_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14944__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ net1262 vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _06501_ _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _07732_ _07735_ _07736_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__o21bai_1
X_10523_ _06087_ net1562 net1023 vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
Xinput19 DAT_I[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11794__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14291_ net1746 _03458_ _03460_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_94_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13242_ net58 _06146_ _06152_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__and3_4
X_16030_ clknet_leaf_157_wb_clk_i _01699_ _00259_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09249__S net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__inv_2
XANTENNA_input73_A wbs_dat_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12183__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15775__A net1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13940__B1 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13173_ _07609_ net382 net293 net1874 vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a22o_1
X_10385_ _03500_ net1076 _05970_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12124_ _04782_ _05280_ net822 vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__or3_1
X_16932_ clknet_leaf_167_wb_clk_i _02601_ _01161_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[905\]
+ sky130_fd_sc_hd__dfrtp_1
X_12055_ _07443_ _07444_ net684 vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__and3_1
X_11006_ _03697_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__xnor2_1
X_16863_ clknet_leaf_157_wb_clk_i _02532_ _01092_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\]
+ sky130_fd_sc_hd__dfrtp_1
X_15814_ clknet_leaf_77_wb_clk_i _01491_ _00041_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16794_ clknet_leaf_33_wb_clk_i _02463_ _01023_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[767\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_412 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15745_ net1294 vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__inv_2
X_12957_ _07247_ net604 net470 net315 net1685 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_29_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13234__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Left_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_104_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11908_ _03632_ _05928_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_138_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15676_ net1281 vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _07588_ net349 net391 net2624 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627_ net1182 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11839_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07317_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__A net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14558_ net1184 vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13509_ _02886_ _02897_ _02899_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a21o_1
X_17277_ team_04_WB.instance_to_wrap.final_design.v_out vssd1 vssd1 vccd1 vccd1 net175
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14489_ net1159 vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09159__S net921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16228_ clknet_leaf_169_wb_clk_i _01897_ _00457_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[201\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13931__B1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16159_ clknet_leaf_154_wb_clk_i _01828_ _00388_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08998__S net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09683__A net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[238\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[206\]
+ net967 vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__mux2_1
XANTENNA__09038__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__A _06932_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ net1101 net1098 vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nor2_1
XANTENNA__12498__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09589__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_143_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09602_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[739\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[707\]
+ net952 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09622__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[261\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09666__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15921__Q net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[934\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[902\]
+ net888 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__mux2_1
XANTENNA__12670__A0 _07356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__S net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09761__S1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__B net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ _04022_ _04023_ _04024_ _04025_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04026_
+ sky130_fd_sc_hd__mux4_1
X_17297__1353 vssd1 vssd1 vccd1 vccd1 _17297__1353/HI net1353 sky130_fd_sc_hd__conb_1
X_09395_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout525_A _06197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_848 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08346_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[474\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__mux2_1
XANTENNA__09513__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__B1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12973__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ _03884_ _03885_ _03886_ _03887_ net788 net809 vssd1 vssd1 vccd1 vccd1 _03888_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12284__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout894_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13922__B1 net104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_142_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09864__Y _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_182_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10170_ _05548_ _05655_ net622 vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__o21a_1
XANTENNA__08701__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11187__X _06676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1106 net1107 vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_4
Xfanout1117 net1118 vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
XANTENNA__12489__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13686__C1 _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1131 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_4
Xfanout1139 net1141 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13860_ net1039 _03247_ _03248_ net1066 net1526 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_87_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09532__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ net254 net2535 net323 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__mux2_1
X_13791_ _03179_ _03180_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12661__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15530_ net1105 vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12742_ _07467_ net348 net403 net2637 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15461_ net1109 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__inv_2
X_12673_ net243 net2537 net475 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__mux2_1
XANTENNA__13205__A2 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14674__A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ clknet_leaf_81_wb_clk_i team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[0\]
+ _01429_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14412_ net1274 vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ net563 _06273_ _06612_ _07105_ _07112_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__a311o_1
XANTENNA__09768__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15392_ net1212 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17131_ clknet_leaf_75_wb_clk_i _02766_ _01360_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_14343_ net1183 vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__inv_2
X_11555_ net532 _06568_ _06572_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10975__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ team_04_WB.instance_to_wrap.CPU_DAT_O\[31\] net1094 net1053 vssd1 vssd1 vccd1
+ vccd1 _06076_ sky130_fd_sc_hd__and3_1
X_17062_ clknet_leaf_49_wb_clk_i _00009_ _01291_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_14274_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[19\] _03448_
+ net819 vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_150_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input76_X net76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _06973_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09268__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire597 team_04_WB.instance_to_wrap.final_design.cpu.Error vssd1 vssd1 vccd1 vccd1
+ net597 sky130_fd_sc_hd__buf_1
XANTENNA__13913__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ net76 team_04_WB.MEM_SIZE_REG_REG\[16\] net982 vssd1 vssd1 vccd1 vccd1 _01678_
+ sky130_fd_sc_hd__mux2_1
X_16013_ clknet_leaf_43_wb_clk_i _01689_ _00242_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12716__B2 _07403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10437_ _06014_ _06015_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09707__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_59_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12192__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _07592_ net373 net291 net1822 vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10368_ _05623_ _05954_ _05955_ net623 net279 vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__o221a_1
XANTENNA__13229__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12107_ net2188 net355 _07508_ net458 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__a22o_1
XANTENNA__12133__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ net228 net2574 net304 vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10299_ _05534_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__or2_1
X_16915_ clknet_leaf_181_wb_clk_i _02584_ _01144_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\]
+ sky130_fd_sc_hd__dfrtp_1
X_12038_ net2276 net515 _07472_ net442 vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XANTENNA__11825__X _07305_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16846_ clknet_leaf_42_wb_clk_i _02515_ _01075_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09442__S net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10588__S net1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16777_ clknet_leaf_122_wb_clk_i _02446_ _01006_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[750\]
+ sky130_fd_sc_hd__dfrtp_1
X_13989_ net1512 net1070 _03329_ net264 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a22o_1
XANTENNA__11273__A team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ net1292 vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__inv_2
XANTENNA__12652__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13995__A3 _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12088__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15659_ net1174 vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08200_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[381\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[299\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[267\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08131_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[702\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[670\]
+ net875 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__mux2_1
X_17329_ net1385 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XFILLER_0_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_170_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10617__A _06140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10966__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08062_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[24\] net1009
+ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__C1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09617__S net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B2 net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__S1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11930__A2 _07008_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[943\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[911\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
X_07915_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__or2_1
XANTENNA__11167__B _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[400\]
+ net873 vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_1
XANTENNA__09431__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout475_A _07662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12891__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09352__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09516_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[804\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\]
+ net882 vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12643__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _03723_ _03947_ _03630_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout907_A net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09378_ _04985_ _04986_ _04987_ _04988_ net791 net802 vssd1 vssd1 vccd1 vccd1 _04989_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08329_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[570\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[538\]
+ net931 vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10527__A team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11340_ net560 _06793_ net573 vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout897_X net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ _06510_ _06759_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_160_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08378__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ net601 _07470_ net469 net310 net1785 vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a32o_1
X_10222_ _05559_ _05647_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__nand2_1
XANTENNA__12174__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10153_ _05686_ _05687_ _05763_ _05684_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_89_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13844__Y _03235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _04502_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\] vssd1
+ vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__and2b_1
X_14961_ net1268 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\] vssd1 vssd1 vccd1
+ vccd1 net1445 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ clknet_leaf_127_wb_clk_i _02369_ _00929_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\]
+ sky130_fd_sc_hd__dfrtp_1
X_13912_ _02982_ _03279_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12882__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14892_ net1119 vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16631_ clknet_leaf_154_wb_clk_i _02300_ _00860_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\]
+ sky130_fd_sc_hd__dfrtp_1
X_13843_ team_04_WB.MEM_SIZE_REG_REG\[31\] _02842_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12189__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12634__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ clknet_leaf_18_wb_clk_i _02231_ _00791_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[535\]
+ sky130_fd_sc_hd__dfrtp_1
X_13774_ net992 _03162_ _03164_ net990 vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__o22a_1
X_10986_ _06346_ _06350_ _06354_ _06474_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and4_1
XFILLER_0_168_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15513_ net1248 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__inv_2
X_12725_ _07450_ net334 net401 net2352 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16493_ clknet_leaf_41_wb_clk_i _02162_ _00722_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15444_ net1235 vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10660__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12656_ net214 net2222 net477 vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
XANTENNA__08606__S net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10708__Y _06197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11607_ net588 net579 net547 vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__mux2_1
X_15375_ net1199 vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__inv_2
XANTENNA__12128__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12587_ net700 _06198_ _07555_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17114_ clknet_leaf_104_wb_clk_i _02749_ _01343_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08161__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14326_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[7\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[6\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[5\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[4\] net1090
+ net1089 vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11538_ _06423_ _07026_ net465 vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__o21ai_1
Xhold408 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\] vssd1 vssd1
+ vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\] vssd1 vssd1
+ vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ clknet_leaf_35_wb_clk_i _02714_ _01274_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
X_14257_ _03438_ _03439_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11469_ _06373_ _06864_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_78_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_748 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13208_ net61 _06145_ _06153_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08341__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188_ _03373_ _03399_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[8\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__11373__B1 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17296__1352 vssd1 vssd1 vccd1 vccd1 _17296__1352/HI net1352 sky130_fd_sc_hd__conb_1
XFILLER_0_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13139_ _07573_ net377 net296 net2055 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_75 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09961__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1108 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[832\] vssd1 vssd1
+ vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[159\] vssd1 vssd1
+ vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12798__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14579__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_10 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11676__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[949\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[917\]
+ net840 vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__B2 net287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12873__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16829_ clknet_leaf_126_wb_clk_i _02498_ _01058_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12625__B1 net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[617\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11979__A2 _07115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_448 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09232_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[490\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[458\]
+ net847 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10651__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09163_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[683\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[651\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13050__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__B1 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08114_ net759 _03622_ _03635_ _03637_ _03644_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o41a_4
X_09094_ net776 _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08045_ _03650_ _03652_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__nor2_4
XFILLER_0_142_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14106__X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold920 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[965\] vssd1 vssd1
+ vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold931 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[76\] vssd1 vssd1
+ vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold942 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\] vssd1 vssd1
+ vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold953 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\] vssd1 vssd1
+ vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[919\] vssd1 vssd1
+ vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09652__S0 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold975 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[77\] vssd1 vssd1
+ vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_A _04166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold986 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\] vssd1 vssd1
+ vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\] vssd1 vssd1
+ vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ net579 _05224_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07943__X _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08947_ _03554_ net703 _04330_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09404__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout857_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11465__X _06954_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12864__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ net778 _04488_ net761 vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14001__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ _03974_ _06306_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12616__B1 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__X _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13959__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09810__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _03696_ net364 _06256_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11641__A net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12510_ _07507_ net482 net424 net2069 vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a22o_1
X_13490_ _03495_ _05808_ net1099 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ net521 net603 _07450_ net428 net1928 vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a32o_1
XANTENNA__13041__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12395__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ _07327_ net2632 net496 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__mux2_1
X_15160_ net1203 vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14111_ team_04_WB.MEM_SIZE_REG_REG\[10\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[10\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__o221a_2
X_11323_ _04247_ net357 vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15091_ net1244 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14042_ net15 net1062 net1038 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1
+ vccd1 vccd1 _01544_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11254_ net566 _06742_ _06739_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12191__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10205_ _05556_ _05650_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11450__S0 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ _06246_ _06578_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10136_ _05717_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__nor2_1
X_15993_ clknet_leaf_71_wb_clk_i _01669_ _00222_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_145_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _04057_ vssd1
+ vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__nor2_1
X_14944_ net1220 vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__inv_2
XANTENNA__12855__B1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11535__B _07023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_141_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14875_ net1145 vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload1_A clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16614_ clknet_leaf_22_wb_clk_i _02283_ _00843_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[587\]
+ sky130_fd_sc_hd__dfrtp_1
X_13826_ net996 _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__nand2_1
XANTENNA__12607__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09720__S net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ clknet_leaf_134_wb_clk_i _02214_ _00774_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09499__Y _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13757_ _02993_ _03098_ _03143_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o31a_1
XANTENNA__13280__B1 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12083__B2 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ _04328_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__nand2_1
XANTENNA__15023__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12708_ net1938 net406 net350 _07357_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11830__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08336__S net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16476_ clknet_leaf_127_wb_clk_i _02145_ _00705_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\]
+ sky130_fd_sc_hd__dfrtp_1
X_13688_ team_04_WB.ADDR_START_VAL_REG\[0\] _03078_ vssd1 vssd1 vccd1 vccd1 _03079_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11830__B2 _04274_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ net1182 vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__inv_2
XANTENNA__13032__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ _07610_ net488 net411 net1657 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08134__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09956__A net639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13583__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ net1215 vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14309_ net178 net68 net101 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__and3b_1
XANTENNA__13478__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold205 net161 vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14073__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15289_ net1245 vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__inv_2
Xhold216 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[560\] vssd1 vssd1
+ vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 net120 vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold238 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\] vssd1 vssd1
+ vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09167__S net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\] vssd1 vssd1
+ vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ clknet_leaf_171_wb_clk_i _02697_ _01257_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08071__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11897__A1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__buf_2
X_09850_ net698 _05451_ _03621_ net905 vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and4b_1
XANTENNA__08211__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout718 net719 vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_6
Xfanout729 net732 vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_165_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_165_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _04387_ _04411_ net662 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__mux2_4
XANTENNA__13099__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net780 _05391_ net763 vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08732_ net729 _04342_ net713 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__o21a_1
XANTENNA__12846__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12310__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ net751 _03662_ _03725_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08594_ net779 _04204_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13271__A0 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout340_A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13810__A2 _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout438_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08246__S net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12276__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09215_ net779 _04825_ net761 vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09146_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[171\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09077_ _04684_ _04685_ _04686_ _04687_ net826 net734 vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10805__A _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_49_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08028_ _03615_ _03623_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and4b_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold750 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[278\] vssd1 vssd1
+ vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10524__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout974_A _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold761 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\] vssd1 vssd1
+ vccd1 vccd1 net2198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold772 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[78\] vssd1 vssd1
+ vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[344\] vssd1 vssd1
+ vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11888__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold794 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[811\] vssd1 vssd1
+ vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09805__S net890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net631 _04839_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12837__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ net604 _07450_ net470 net311 net1886 vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__a32o_1
XANTENNA__14012__A _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11941_ _03631_ _05967_ net696 _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__a211o_1
XFILLER_0_169_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08600__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16000__Q team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14660_ net1169 vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__inv_2
X_11872_ team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] _07236_ _07345_ _07239_ vssd1
+ vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__a31o_1
XFILLER_0_169_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09540__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13611_ _02997_ net1077 _07693_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__or4bb_1
X_10823_ _03753_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_49_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14591_ net1182 vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__inv_2
XANTENNA__12065__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13062__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ clknet_leaf_110_wb_clk_i _01999_ _00559_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\]
+ sky130_fd_sc_hd__dfrtp_1
X_13542_ _02930_ _02931_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__or2_1
XANTENNA__11812__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10754_ net640 net543 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__and2_1
X_17295__1351 vssd1 vssd1 vccd1 vccd1 _17295__1351/HI net1351 sky130_fd_sc_hd__conb_1
XFILLER_0_94_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16261_ clknet_leaf_6_wb_clk_i _01930_ _00490_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13473_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__inv_2
X_10685_ net2591 net711 _06180_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a22o_1
XANTENNA__13014__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15212_ net1121 vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__inv_2
X_12424_ net525 net610 _07397_ net435 net1567 vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_97_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16192_ clknet_leaf_141_wb_clk_i _01861_ _00421_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15143_ net1139 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ net228 net670 vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__and2_2
XFILLER_0_106_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11306_ _06575_ _06580_ net539 vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__mux2_1
X_12286_ net222 net674 vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__and2_1
X_15074_ net1255 vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14025_ _07688_ net1041 _03349_ net1072 net1506 vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a32o_1
X_11237_ _04328_ _04357_ net357 vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__or3_1
XANTENNA__11879__A1 _03613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08744__B2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09715__S net969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_143_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ _06470_ _06474_ _06350_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_143_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13237__S net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] _05223_ vssd1
+ vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12141__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15976_ clknet_leaf_51_wb_clk_i _01652_ _00205_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12828__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11099_ _06582_ _06587_ net560 vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_160_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_160_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14927_ net1140 vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__inv_2
X_14858_ net1112 vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_69_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09450__S net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13809_ _03194_ _03199_ _02948_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__a21oi_1
XANTENNA__14068__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__B2 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14789_ net1111 vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08355__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11803__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ clknet_leaf_192_wb_clk_i _02197_ _00757_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[501\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11803__B2 _04004_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12096__B net679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15688__A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13005__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16459_ clknet_leaf_25_wb_clk_i _02128_ _00688_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[432\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[14\] team_04_WB.instance_to_wrap.CPU_DAT_O\[14\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__mux2_4
XFILLER_0_54_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _04031_ net595 _04084_ _04029_ net640 vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout504 net506 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_8
Xfanout515 _07449_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_6
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout526 _06195_ vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_6
XANTENNA__11727__Y _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09833_ _04611_ _04669_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout537 net538 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__clkbuf_4
Xfanout548 _05377_ vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__buf_2
XANTENNA__09852__C _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout559 _05309_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout388_A _07673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ net719 _05367_ _05373_ _05361_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__a31o_4
XFILLER_0_77_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_167_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_167_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08715_ _04322_ _04323_ _04324_ _04325_ net787 net810 vssd1 vssd1 vccd1 vccd1 _04326_
+ sky130_fd_sc_hd__mux4_1
X_09695_ _05300_ _05305_ net724 vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout555_A net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_A net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08646_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[149\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09360__S net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08577_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[758\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__mux2_1
XANTENNA__12598__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_475 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1252_X net1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] _06039_
+ _06041_ _06033_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08649__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13011__A3 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ net730 _04733_ net714 vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_40_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12140_ _07333_ net2619 net512 vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XANTENNA__12770__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12071_ net2068 net353 _07490_ net445 vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[296\] vssd1 vssd1
+ vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[639\] vssd1 vssd1
+ vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ team_04_WB.MEM_SIZE_REG_REG\[19\] _06510_ vssd1 vssd1 vccd1 vccd1 _06511_
+ sky130_fd_sc_hd__or2_2
XANTENNA__09535__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13057__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15830_ clknet_leaf_93_wb_clk_i _01507_ _00057_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13852__Y _03243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15761_ net1275 vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__inv_2
XANTENNA__13483__B1 team_04_WB.ADDR_START_VAL_REG\[28\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ net610 _07357_ net474 net317 net1569 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__a32o_1
XANTENNA__08946__Y _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14712_ net1203 vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__inv_2
X_11924_ net651 net251 vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15692_ net1268 vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__inv_2
XANTENNA__14027__A2 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13235__A0 net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14643_ net1227 vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07331_ sky130_fd_sc_hd__a21o_1
XANTENNA__12038__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12197__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12589__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _06286_ _06293_ _05463_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_99_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14574_ net1263 vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__inv_2
XANTENNA__13786__B2 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11786_ net652 net219 vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08888__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16313_ clknet_leaf_177_wb_clk_i _01982_ _00542_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[286\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ net989 _02915_ _02913_ net994 vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17293_ net1349 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10737_ net564 net546 net540 vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_136_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16244_ clknet_leaf_4_wb_clk_i _01913_ _00473_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[217\]
+ sky130_fd_sc_hd__dfrtp_1
X_13456_ net992 _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10668_ net1570 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1
+ vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a22o_1
XANTENNA__13002__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12407_ net2174 net432 _07631_ net520 vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_114_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12136__S net511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16175_ clknet_leaf_3_wb_clk_i _01844_ _00404_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\]
+ sky130_fd_sc_hd__dfrtp_1
X_13387_ _07809_ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__and2_1
X_10599_ team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] net1096 net1051 vssd1 vssd1 vccd1
+ vccd1 _06138_ sky130_fd_sc_hd__and3_1
XANTENNA__12210__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09793__X _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput118 net118 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__clkbuf_4
X_15126_ net1221 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__inv_2
XANTENNA__12761__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput129 net129 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__clkbuf_4
X_12338_ net2371 net499 _07613_ net437 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15057_ net1266 vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__inv_2
X_12269_ net2358 net503 _07577_ net439 vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a22o_1
XANTENNA__09065__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08717__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ _05137_ net264 _03335_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_162_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_133_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15959_ clknet_4_13__leaf_wb_clk_i _01635_ _00188_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13474__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12277__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A1 _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _04105_ _04110_ net770 vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09480_ _05087_ _05088_ _05089_ _05090_ net792 net802 vssd1 vssd1 vccd1 vccd1 _05091_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09180__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08431_ _04038_ _04039_ _04040_ _04041_ net785 net800 vssd1 vssd1 vccd1 vccd1 _04042_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08362_ _03960_ _03961_ _03972_ net717 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a22o_2
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08293_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[27\]
+ net860 vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08405__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_172_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout303_A _07681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1045_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12752__A2 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11960__B1 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14114__X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout301 _07682_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_4
XANTENNA__12504__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09355__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout323 _07671_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_4
Xfanout334 net336 vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout672_A _07554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 net351 vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_4
X_17294__1350 vssd1 vssd1 vccd1 vccd1 _17294__1350/HI net1350 sky130_fd_sc_hd__conb_1
Xfanout367 net372 vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__buf_4
X_09816_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[769\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__mux2_1
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_4
Xfanout389 _07673_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_4
XFILLER_0_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10521__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\]
+ net903 vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09678_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[354\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[322\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09090__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12448__C net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ net465 _07120_ net285 vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11779__B1 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11571_ team_04_WB.MEM_SIZE_REG_REG\[5\] _06500_ vssd1 vssd1 vccd1 vccd1 _07060_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11243__A2 _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13310_ net1083 team_04_WB.MEM_SIZE_REG_REG\[23\] vssd1 vssd1 vccd1 vccd1 _07736_
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_162_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10522_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[26\]
+ _06086_ net1050 vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__mux2_1
XANTENNA__12991__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14290_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[25\] _03458_
+ net818 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08434__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09819__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10453_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _06028_
+ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__xor2_1
X_13241_ net69 team_04_WB.MEM_SIZE_REG_REG\[0\] net985 vssd1 vssd1 vccd1 vccd1 _01662_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08947__A1 _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12743__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input66_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ net282 _05968_ _05969_ _05966_ net1057 vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a221o_1
X_13172_ _07608_ net383 net292 net1740 vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12123_ net2048 net355 _07516_ net460 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
XANTENNA__12480__A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09265__S net925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12054_ net2580 net517 _07480_ net457 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a22o_1
X_16931_ clknet_leaf_122_wb_clk_i _02600_ _01160_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08022__X _03633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11096__A _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _03753_ _05463_ _06311_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__o21ba_1
X_16862_ clknet_leaf_129_wb_clk_i _02531_ _01091_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
X_16793_ clknet_leaf_154_wb_clk_i _02462_ _01022_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12259__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15744_ net1293 vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ net699 _06183_ _07666_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_29_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10090__A_N _04612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ team_04_WB.instance_to_wrap.CPU_DAT_O\[11\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07376_ sky130_fd_sc_hd__a21o_1
X_15675_ net1281 vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__inv_2
XANTENNA__11482__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _07587_ net344 net390 net2110 vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10690__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14626_ net1255 vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_103_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ net704 _05862_ _07315_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14557_ net1178 vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_155_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ _06525_ _06591_ net690 vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__a21o_1
XANTENNA__12431__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13508_ _02884_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17276_ net1335 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12982__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08344__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14488_ net1251 vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__inv_2
Xclkbuf_4_0__f_wb_clk_i clknet_3_0_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_130_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16227_ clknet_leaf_121_wb_clk_i _01896_ _00456_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\]
+ sky130_fd_sc_hd__dfrtp_1
X_13439_ _07856_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__nor2_1
XANTENNA__10606__C _06141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13931__A1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09964__A _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12734__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ clknet_leaf_157_wb_clk_i _01827_ _00387_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[131\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15109_ net1108 vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__inv_2
XANTENNA__14081__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ clknet_leaf_177_wb_clk_i _01758_ _00318_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_08980_ _04587_ _04588_ _04589_ _04590_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04591_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09038__S1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07931_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\] net1080
+ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nor2_1
XANTENNA__12498__A1 _07495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09601_ _05208_ _05209_ _05210_ _05211_ net794 net813 vssd1 vssd1 vccd1 vccd1 _05212_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_127_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09532_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[325\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[966\]
+ net888 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout253_A _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10681__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08414_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[697\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\]
+ net839 vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09698__X _05309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09394_ _03724_ _03893_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10069__B _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12422__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08345_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[314\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout420_A _07658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14109__X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1162_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout518_A _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08276_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[699\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[667\]
+ net929 vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12284__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__A1 _04328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout306_X net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13922__B2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12489__A1 _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_182_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_182_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xfanout1107 net1115 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13686__B1 net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1118 net1123 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1129 net1131 vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__buf_2
XANTENNA__14004__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_35_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__S net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12810_ _07374_ net2438 net323 vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13790_ _03180_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__inv_2
XANTENNA__08429__S net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _07466_ net350 net402 net2297 vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08865__B1 _04439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ net1171 vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__inv_2
XANTENNA__10672__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12672_ net255 net2476 net478 vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14411_ net1274 vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _05404_ net533 _06257_ _07106_ net465 vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__a311o_1
X_15391_ net1273 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__inv_2
XANTENNA__12413__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13610__B1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ clknet_leaf_75_wb_clk_i net1516 _01359_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_133_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14342_ net1183 vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12964__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08164__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ _05336_ net547 net532 _06569_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a211o_1
X_17061_ clknet_leaf_49_wb_clk_i _00008_ _01290_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10505_ _05999_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14273_ _03448_ _03449_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ team_04_WB.MEM_SIZE_REG_REG\[12\] _06505_ vssd1 vssd1 vccd1 vccd1 _06974_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_150_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14690__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09268__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16012_ clknet_leaf_51_wb_clk_i _01688_ _00241_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_13224_ net77 team_04_WB.MEM_SIZE_REG_REG\[17\] net985 vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12716__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10436_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06013_
+ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and2_1
XANTENNA_input69_X net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13155_ net699 _07590_ _07666_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__or3_4
X_10367_ _05745_ _05747_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__xnor2_1
X_12106_ net249 net679 vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__and2_1
X_10298_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[15\] _05533_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a21oi_1
X_13086_ net221 net2562 net305 vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13141__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ net251 net680 vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__and2_1
X_16914_ clknet_leaf_9_wb_clk_i _02583_ _01143_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16845_ clknet_leaf_42_wb_clk_i _02514_ _01074_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[818\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13245__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16776_ clknet_leaf_160_wb_clk_i _02445_ _01005_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13988_ _04752_ _03326_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__nor2_1
XANTENNA__08339__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12101__B1 _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ net1294 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_137_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12939_ net259 net2142 net319 vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14865__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10663__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15658_ net1174 vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__inv_2
XANTENNA__09959__A _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08863__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ net1267 vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08608__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14076__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15589_ net1108 vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__inv_2
XANTENNA__10415__A0 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08130_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[766\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[734\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__mux2_1
X_17328_ net1384 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__09030__Y _04641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08074__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10966__A1 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ net722 _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__or2_1
X_17259_ net1319 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_4_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12707__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1007\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[975\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_07914_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__nor2_1
XANTENNA__13132__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\]
+ net873 vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
XANTENNA__09431__S1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__B1 _07614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__A team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09860__C net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09639__A2 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13950__Y _03309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[868\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\]
+ net881 vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__mux2_1
XANTENNA__12643__A1 _07614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout635_A _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ net626 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[7\]
+ net945 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout802_A net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12295__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_348 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1165_X net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08328_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[634\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10527__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ team_04_WB.MEM_SIZE_REG_REG\[17\] _06509_ team_04_WB.MEM_SIZE_REG_REG\[18\]
+ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08712__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__B1 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] net1055 _05822_
+ _05825_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10152_ _05688_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16003__Q team_04_WB.MEM_SIZE_REG_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _04441_ vssd1
+ vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__or2_1
X_14960_ net1163 vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11134__A1 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[30\]
+ vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09878__A2 _04610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ _03281_ _03284_ net2099 net1067 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_input29_A DAT_I[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ net1160 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__inv_2
XANTENNA__13065__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ clknet_leaf_14_wb_clk_i _02299_ _00859_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\]
+ sky130_fd_sc_hd__dfrtp_1
X_13842_ _07876_ _02845_ _02844_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16561_ clknet_leaf_176_wb_clk_i _02230_ _00790_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13773_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _05879_ net1099
+ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__mux2_1
XANTENNA__12634__A1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10985_ _06459_ _06462_ _06472_ _06473_ _06458_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__a32o_1
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14685__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12757__X _07670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15512_ net1205 vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__inv_2
X_12724_ net701 _07448_ _07663_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__or3_4
X_16492_ clknet_leaf_107_wb_clk_i _02161_ _00721_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ net1233 vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ net212 net2466 net477 vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
XANTENNA__10718__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_152_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11606_ _07094_ _05473_ _07093_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__or3b_1
XFILLER_0_167_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15374_ net1207 vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12586_ _07553_ net494 net419 net1745 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14139__A1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17113_ clknet_leaf_104_wb_clk_i _02748_ _01342_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14325_ _03476_ _03482_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08161__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ _06396_ _06422_ _06392_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold409 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\] vssd1 vssd1
+ vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
X_17044_ clknet_leaf_1_wb_clk_i _02713_ _01273_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
X_14256_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\] _03437_
+ net820 vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11468_ net755 _06915_ _06917_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08622__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13207_ net61 _06145_ _06153_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__and3_4
XANTENNA__09110__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _03532_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__o21ai_1
X_14187_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] _03368_
+ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
XANTENNA__12144__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11373__A1 team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10176__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _04754_ net365 vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nor2_1
XANTENNA__12570__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _07572_ net374 net295 net1929 vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13764__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13069_ net260 net2491 net303 vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__mux2_1
Xhold1109 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\] vssd1 vssd1
+ vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12322__B1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16828_ clknet_leaf_125_wb_clk_i _02497_ _01057_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16759_ clknet_leaf_155_wb_clk_i _02428_ _00988_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _04907_ _04908_ _04909_ _04910_ net826 net742 vssd1 vssd1 vccd1 vccd1 _04911_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09231_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[298\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[266\]
+ net848 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12389__A0 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08057__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09162_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[715\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08113_ _03637_ _03722_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__or2_2
X_09093_ _04700_ _04701_ _04702_ _04703_ net796 net816 vssd1 vssd1 vccd1 vccd1 _04704_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13737__A1_N net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_839 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09628__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__B1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08044_ net1078 net1030 net1026 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__o31a_2
XANTENNA__08532__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold910 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\] vssd1 vssd1
+ vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[843\] vssd1 vssd1
+ vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11349__D1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold932 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[913\] vssd1 vssd1
+ vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[974\] vssd1 vssd1
+ vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11459__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold954 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\] vssd1 vssd1
+ vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold965 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\] vssd1 vssd1
+ vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__A1 _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[157\] vssd1 vssd1
+ vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09652__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold987 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\] vssd1 vssd1
+ vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[924\] vssd1 vssd1
+ vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ net579 _05224_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout585_A net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_134_Left_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13105__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _04556_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__inv_2
XANTENNA__14122__X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09404__S1 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _04484_ _04485_ _04486_ _04487_ net789 net801 vssd1 vssd1 vccd1 vccd1 _04488_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11824__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10770_ net645 _03695_ net357 vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__or3_1
XANTENNA__08707__S net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_143_Left_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11641__B _07129_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[230\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12456__C net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12919__A2 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ net699 _06198_ _07448_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__or3_4
XFILLER_0_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13592__A2 net271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net246 net2558 net495 vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ team_04_WB.MEM_SIZE_REG_REG\[9\] net987 net980 team_04_WB.ADDR_START_VAL_REG\[9\]
+ net1004 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__o221a_2
XANTENNA__09538__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _06790_ _06800_ _06810_ net288 vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__a22o_1
X_15090_ net1245 vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__inv_2
XANTENNA__11369__A net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ net16 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1
+ vccd1 vccd1 _01545_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_56_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11253_ net553 _06663_ _06740_ _06531_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_127_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_152_Left_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10204_ _05674_ _05769_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11184_ _04194_ net363 _06670_ _06672_ net287 vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_73_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10135_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _04948_ vssd1
+ vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15992_ clknet_leaf_71_wb_clk_i _01668_ _00221_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_145_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10066_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _04057_ vssd1
+ vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__and2_1
X_14943_ net1270 vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_174_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11658__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ net1151 vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13825_ net989 _03215_ _03213_ net994 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a2bb2o_1
X_16613_ clknet_leaf_170_wb_clk_i _02282_ _00842_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[586\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12487__X _07656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_161_Left_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16544_ clknet_leaf_139_wb_clk_i _02213_ _00773_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[517\]
+ sky130_fd_sc_hd__dfrtp_1
X_13756_ _02957_ _02966_ _02970_ _03146_ _02956_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__o221a_1
XFILLER_0_174_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13280__A1 _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ _04357_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__xor2_2
XANTENNA__12083__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11551__B _07039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ net1999 net404 net338 _07350_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16475_ clknet_leaf_101_wb_clk_i _02144_ _00704_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[448\]
+ sky130_fd_sc_hd__dfrtp_1
X_13687_ net710 _03075_ _03076_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__o22a_1
XANTENNA__12139__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10899_ net659 _06284_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__nor2_1
X_15426_ net1239 vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__inv_2
XANTENNA__08039__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13032__A1 _07493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12638_ _07609_ net492 net411 net1737 vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08134__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13583__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ net1149 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _07536_ net493 net418 net1707 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12791__A0 net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14308_ _03621_ net754 _04784_ net691 vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.Error
+ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_117_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15288_ net1205 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__inv_2
Xhold206 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[118\] vssd1 vssd1
+ vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08352__S net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold217 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[189\] vssd1 vssd1
+ vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\] vssd1 vssd1
+ vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_170_Left_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17027_ clknet_leaf_122_wb_clk_i _02696_ _01256_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_169_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold239 net129 vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
X_14239_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[6\] _03426_ vssd1
+ vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_169_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10149__A2 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08211__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 _03627_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout719 _03674_ vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_165_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ net717 _04410_ _04399_ _04398_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__o2bb2a_2
X_09780_ _05387_ _05388_ _05389_ _05390_ net794 net802 vssd1 vssd1 vccd1 vccd1 _05391_
+ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10911__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08731_ _04338_ _04339_ _04340_ _04341_ net829 net735 vssd1 vssd1 vccd1 vccd1 _04342_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_63 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1290 net1293 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_89_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08662_ net766 _04272_ _04261_ _04255_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o2bb2a_4
X_08593_ _04200_ _04201_ _04202_ _04203_ net783 net800 vssd1 vssd1 vccd1 vccd1 _04204_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15811__30 clknet_leaf_62_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__inv_2
XANTENNA__11806__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13810__A3 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout333_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _04821_ _04822_ _04823_ _04824_ net784 net800 vssd1 vssd1 vccd1 vccd1 _04825_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[235\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[203\]
+ net915 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__mux2_1
XANTENNA__10645__X _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout500_A _07591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1242_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12782__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09358__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09076_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[556\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[524\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__mux2_1
XANTENNA__08115__X _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12292__B _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _03617_ _03597_ _03609_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__or3b_1
XANTENNA__13956__X _03312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\] vssd1 vssd1
+ vccd1 vccd1 net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\] vssd1 vssd1
+ vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10524__C net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold762 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\] vssd1 vssd1
+ vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold773 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\] vssd1 vssd1
+ vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[506\] vssd1 vssd1
+ vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[597\] vssd1 vssd1
+ vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_89_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_09978_ net633 _04787_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_08929_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11940_ net756 _05968_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ _05466_ _07240_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__or2_2
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ net1102 _05959_ net995 _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10822_ _03861_ _06310_ net657 vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__o21a_1
XANTENNA__13262__A1 team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14590_ net1184 vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__inv_2
XANTENNA__12065__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__X _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13541_ _02931_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__inv_2
XANTENNA__09561__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10753_ _03892_ _03946_ net550 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16260_ clknet_leaf_169_wb_clk_i _01929_ _00489_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[233\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _02856_ _02862_ team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1
+ _02863_ sky130_fd_sc_hd__a21oi_1
XANTENNA_input96_A wbs_dat_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\] _06179_ _06180_
+ net34 vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15211_ net1161 vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__inv_2
X_12423_ net520 net602 _07391_ net432 net1603 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_164_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16191_ clknet_leaf_155_wb_clk_i _01860_ _00420_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12773__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15142_ net1104 vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__inv_2
XFILLER_0_65_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12354_ net2234 net501 _07621_ net455 vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _06792_ _06793_ net560 vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__mux2_1
X_15073_ net1188 vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__inv_2
XFILLER_0_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ net2536 net505 _07585_ net456 vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a22o_1
X_14024_ _07694_ _03348_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_147_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11236_ _06279_ _06724_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_112_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08900__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_123_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ net706 _06651_ _06654_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_143_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[3\] _05223_ vssd1
+ vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__and2_1
X_15975_ clknet_leaf_50_wb_clk_i _01651_ _00204_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11098_ _06584_ _06586_ net537 vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_160_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10049_ _03591_ _04784_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__or2_1
X_14926_ net1198 vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14857_ net1136 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13253__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11562__A _05336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13808_ _02947_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__and2b_1
XANTENNA__12056__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08347__S net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14788_ net1168 vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13739_ team_04_WB.ADDR_START_VAL_REG\[9\] _03123_ _03126_ _03129_ vssd1 vssd1 vccd1
+ vccd1 _03130_ sky130_fd_sc_hd__and4_1
X_16527_ clknet_leaf_187_wb_clk_i _02196_ _00756_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08355__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09967__A _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13005__A1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16458_ clknet_leaf_163_wb_clk_i _02127_ _00687_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14202__B1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15409_ net1276 vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__inv_2
XANTENNA__14084__S net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16389_ clknet_leaf_170_wb_clk_i _02058_ _00618_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10906__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12764__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_162_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09178__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08432__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12516__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _03920_ net642 _03975_ _03919_ _03891_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__a32o_1
XANTENNA__08810__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 net506 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__clkbuf_8
Xfanout516 _07449_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_4
XFILLER_0_158_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09832_ _04611_ _04725_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__or2_1
Xfanout527 _06195_ vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_171_Right_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout538 _05434_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09852__D net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_2
X_09763_ net719 _05367_ _05373_ _05361_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__a31oi_4
XANTENNA__08111__A net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
X_09694_ _05301_ _05302_ _05303_ _05304_ net834 net746 vssd1 vssd1 vccd1 vccd1 _05305_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_174_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08645_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__mux2_1
XANTENNA__09791__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout450_A net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[534\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_136_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_X net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12755__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09128_ net726 _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12507__B1 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09816__S net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12070_ net227 net677 vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__and2_2
Xhold570 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\] vssd1 vssd1
+ vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[185\] vssd1 vssd1
+ vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\] vssd1 vssd1
+ vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ team_04_WB.MEM_SIZE_REG_REG\[18\] team_04_WB.MEM_SIZE_REG_REG\[17\] _06509_
+ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__or3_1
XANTENNA__13180__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15119__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__A team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11730__A1 _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15760_ net1290 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__inv_2
X_12972_ net605 _07350_ net470 net314 net1560 vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a32o_1
XANTENNA__10297__A1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A DAT_I[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ net695 _06991_ _07389_ net615 vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__a211oi_1
X_14711_ net1228 vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__inv_2
X_15691_ net1256 vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__inv_2
XANTENNA__11494__B1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15850__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12478__A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13073__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14642_ net1237 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__inv_2
X_11854_ net704 _05875_ _07329_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12038__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__B net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ _05463_ _06293_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__or2_1
X_14573_ net1264 vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11785_ net613 _07269_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__and3_2
XFILLER_0_131_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13524_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\] _05845_ net1099
+ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__mux2_1
X_16312_ clknet_leaf_152_wb_clk_i _01981_ _00541_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[285\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12994__B1 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17292_ net1348 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10736_ _06217_ _06224_ net574 vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__mux2_1
XANTENNA_input99_X net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08691__A _04273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16243_ clknet_leaf_185_wb_clk_i _01912_ _00472_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[216\]
+ sky130_fd_sc_hd__dfrtp_1
X_13455_ _07876_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__xor2_2
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ net1546 net1019 net1015 team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1
+ vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12746__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ net651 net601 net240 vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16174_ clknet_leaf_29_wb_clk_i _01843_ _00403_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\]
+ sky130_fd_sc_hd__dfrtp_1
X_13386_ _07805_ _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__or2_1
XANTENNA__12210__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ _06137_ net1860 net1022 vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15125_ net1209 vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ net253 net668 vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__and2_1
Xoutput119 net119 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__clkbuf_4
X_15056_ net1164 vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_110_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ net254 net672 vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__and2_1
XANTENNA__13248__S net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ net1538 net1069 _03339_ net264 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__a22o_1
XANTENNA__13171__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15029__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ net464 _06688_ _06701_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_162_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12152__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__A0 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ net243 net647 vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__and2_1
XANTENNA__14120__C1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15958_ clknet_leaf_79_wb_clk_i _01634_ _00187_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12277__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ net1155 vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15889_ clknet_leaf_99_wb_clk_i _01566_ _00116_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08350__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[24\]
+ net917 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17343__1399 vssd1 vssd1 vccd1 vccd1 _17343__1399/HI net1399 sky130_fd_sc_hd__conb_1
XANTENNA__13226__A1 team_04_WB.MEM_SIZE_REG_REG\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08361_ _03966_ _03971_ net722 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11788__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_914 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12985__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09697__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[123\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08805__S net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12737__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08405__A1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07945__A team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09636__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13162__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout498_A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout313 _07678_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout324 net325 vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_6
Xfanout335 net336 vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
Xfanout346 net348 vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
Xfanout357 net359 vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_2
X_09815_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[865\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\]
+ net893 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__mux2_1
XANTENNA_input3_A DAT_I[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout368 net372 vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_2
Xfanout379 net381 vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[160\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__mux2_1
XANTENNA__09371__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ _05284_ _05285_ _05286_ _05287_ net835 net745 vssd1 vssd1 vccd1 vccd1 _05288_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08628_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[756\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[724\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
XANTENNA__13217__A1 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08559_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\]
+ net850 vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12976__B1 net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ team_04_WB.MEM_SIZE_REG_REG\[0\] _07058_ vssd1 vssd1 vccd1 vccd1 _07059_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10521_ team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] net1096 net1053 vssd1 vssd1 vccd1
+ vccd1 _06086_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__B1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09819__S1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ net80 team_04_WB.MEM_SIZE_REG_REG\[1\] net985 vssd1 vssd1 vccd1 vccd1 _01663_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10452_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _06028_
+ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08947__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13171_ _07607_ net375 net291 net1781 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a22o_1
XANTENNA__11400__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13940__A2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383_ net618 _05967_ net282 vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11951__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09546__S net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_12122_ _07443_ _07444_ net679 vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__and3_2
XANTENNA_input59_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12480__B net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13068__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13153__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16930_ clknet_leaf_147_wb_clk_i _02599_ _01159_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[903\]
+ sky130_fd_sc_hd__dfrtp_1
X_12053_ net228 net682 vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__and2_1
XANTENNA__11703__A1 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _06315_ _06318_ _06491_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__and3_1
XANTENNA__12900__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11096__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ clknet_leaf_132_wb_clk_i _02530_ _01090_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14688__A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14102__C1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout880 net883 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__clkbuf_4
Xfanout891 net895 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
X_16792_ clknet_leaf_156_wb_clk_i _02461_ _01021_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12259__A2 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15743_ net1290 vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__inv_2
X_12955_ _07445_ net2598 net321 vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__mux2_1
XANTENNA__09755__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14200__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ net2331 net527 net449 _07375_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15674_ net1183 vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__inv_2
X_12886_ _07586_ net344 net390 net1935 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11837_ net757 _05857_ _06185_ _04219_ net689 vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14625_ net1148 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12967__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17344_ net1400 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
X_14556_ net1184 vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _03631_ _05781_ net694 _07255_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__a211o_1
XANTENNA__12431__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09310__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ _02885_ _02895_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__and2b_1
X_10719_ net586 _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__nor2_1
X_17275_ net1334 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__12147__S net512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14487_ net1119 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11699_ net572 _06745_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__nor2_1
XANTENNA__12719__B1 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ _07729_ _07863_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__nand2_1
X_16226_ clknet_leaf_144_wb_clk_i _01895_ _00455_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13767__A team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11839__X _07317_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ clknet_leaf_130_wb_clk_i _01826_ _00386_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13931__A2 net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\] team_04_WB.MEM_SIZE_REG_REG\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08494__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09456__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ net1171 vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16088_ clknet_leaf_153_wb_clk_i _01757_ _00317_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13144__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\] net1077
+ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__or2_1
X_15039_ net1242 vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__inv_2
XANTENNA__12498__A2 net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09980__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09600_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[931\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[899\]
+ net958 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09531_ _05110_ net587 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__xnor2_1
X_09462_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[806\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[774\]
+ net888 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08413_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[761\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10681__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ net589 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout246_A _07320_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12958__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08344_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[378\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[346\]
+ net861 vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08535__S net917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12422__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11225__A3 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08275_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout413_A net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12973__A3 net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1155_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13135__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1110 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12489__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13686__B2 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1119 net1123 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__buf_4
XFILLER_0_100_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11449__A0 _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09729_ _05337_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__or2_4
Xclkbuf_leaf_151_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_151_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__13989__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ _07465_ net338 net400 net1876 vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08865__A1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10672__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ net257 net2587 net478 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12949__A0 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14410_ net1267 vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__inv_2
XANTENNA__11660__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ net569 _06987_ _06278_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15390_ net1236 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13610__A1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12413__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ net1183 vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _05464_ _06201_ _05469_ _05518_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__or4b_1
XANTENNA__10975__A2 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17060_ clknet_leaf_49_wb_clk_i _00038_ _01289_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10504_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and2b_1
X_14272_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\] _03447_
+ net819 vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__o21ai_1
X_11484_ net708 _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__nor2_1
XFILLER_0_162_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16011_ clknet_leaf_43_wb_clk_i _01687_ _00240_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_13223_ net78 team_04_WB.MEM_SIZE_REG_REG\[18\] net982 vssd1 vssd1 vccd1 vccd1 _01680_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_150_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13913__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06013_
+ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__nor2_1
XANTENNA__13587__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__S net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ _07588_ net382 net297 net2113 vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08180__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ _05595_ _05621_ _05622_ net624 vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__o31ai_1
XANTENNA__08033__X _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342__1398 vssd1 vssd1 vccd1 vccd1 _17342__1398/HI net1398 sky130_fd_sc_hd__conb_1
XANTENNA__13126__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12105_ net2154 net353 _07507_ net441 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__a22o_1
X_13085_ net229 net2387 net304 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__mux2_1
X_10297_ net624 _05892_ net278 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__o21ai_1
X_16913_ clknet_leaf_176_wb_clk_i _02582_ _01142_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\]
+ sky130_fd_sc_hd__dfrtp_1
X_12036_ net2523 net515 _07471_ net439 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11835__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16844_ clknet_leaf_118_wb_clk_i _02513_ _01073_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[817\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16775_ clknet_leaf_21_wb_clk_i _02444_ _01004_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13987_ net1528 net1070 _03328_ net265 vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12101__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15726_ net1296 vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__inv_2
X_12938_ _07340_ net2407 net321 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12652__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ net1174 vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__inv_2
XANTENNA__10663__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__X _06227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ _07569_ net339 net389 net2083 vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_174_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15042__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ net1282 vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_174_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15588_ net1171 vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327_ net1383 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11612__B1 _06948_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539_ net1286 vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__inv_2
XANTENNA__14881__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__A _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ _03664_ _03665_ _03669_ _03670_ net827 net735 vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17258_ net1318 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_153_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16209_ clknet_leaf_172_wb_clk_i _01878_ _00438_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14092__S net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17189_ clknet_leaf_78_wb_clk_i _02801_ _01418_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10179__B1 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10914__A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A1 _03632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__B2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08090__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__Y _05800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[783\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__mux2_1
X_07913_ team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[1\] team_04_WB.instance_to_wrap.final_design.vga.v_current_state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__and2b_1
X_08893_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[304\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\]
+ net873 vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__mux2_1
XANTENNA__07942__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12891__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout363_A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ net730 _05124_ net714 vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_56_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12643__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__B2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09445_ net767 _05055_ _05044_ _05043_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10654__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[27\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout628_A _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09376_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[103\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[71\]
+ net950 vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12295__B net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ net772 _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__or2_1
XANTENNA__11603__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1158_X net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__C net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__A _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[507\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[475\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10824__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08189_ _03796_ _03797_ _03798_ _03799_ net832 net737 vssd1 vssd1 vccd1 vccd1 _03800_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09096__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13200__A _03548_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ net277 _05824_ net1074 vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13108__B1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _05691_ _05760_ _05689_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_37_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _04441_ vssd1
+ vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _02969_ _02980_ _03280_ _03243_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a31o_1
XANTENNA__14031__A team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ net1116 vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__inv_2
XANTENNA__12882__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _06499_ net272 net709 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_211 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13772_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] net1044 _03162_
+ net1081 vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__o22a_1
X_16560_ clknet_leaf_191_wb_clk_i _02229_ _00789_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[533\]
+ sky130_fd_sc_hd__dfrtp_1
X_10984_ _04328_ _06457_ _06461_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12634__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__Y _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15511_ net1233 vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
X_12723_ net2592 net407 net349 _07446_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a22o_1
X_16491_ clknet_leaf_16_wb_clk_i _02160_ _00720_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[464\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13081__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15442_ net1247 vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__inv_2
X_12654_ net211 net2344 net476 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _05252_ _06248_ _06273_ _06632_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__a22o_1
X_15373_ net1201 vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__inv_2
X_12585_ _07552_ net489 net418 net1726 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a22o_1
XANTENNA__08697__S0 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input81_X net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17112_ clknet_leaf_104_wb_clk_i _02747_ _01341_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11536_ team_04_WB.MEM_SIZE_REG_REG\[6\] _06501_ vssd1 vssd1 vccd1 vccd1 _07025_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14324_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[11\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[10\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[9\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[8\] net1091
+ net1089 vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux4_1
XANTENNA__11070__A1 _03946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08471__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14255_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\] _03437_
+ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__and2_1
X_17043_ clknet_leaf_181_wb_clk_i _02712_ _01272_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
X_11467_ _06935_ _06955_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13206_ _03516_ _07699_ net1072 _07702_ team_04_WB.instance_to_wrap.BUSY_O vssd1
+ vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__o32a_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_78_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14186_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ _03372_ _03391_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__and4_1
XANTENNA__11549__B _07037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09110__S1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11398_ net466 _06884_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__nand2_1
X_13137_ _07571_ net382 net297 net2192 vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__a22o_1
X_10349_ _05626_ net623 _05936_ _05938_ net282 vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a311o_1
X_13068_ net246 net2583 net302 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12019_ net245 net681 vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__and2_1
XANTENNA__15037__A net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_79_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12873__A2 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16827_ clknet_leaf_97_wb_clk_i _02496_ _01056_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[800\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16758_ clknet_leaf_15_wb_clk_i _02427_ _00987_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[731\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08829__A1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12625__A2 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15709_ net1281 vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12396__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16689_ clknet_leaf_176_wb_clk_i _02358_ _00918_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10909__A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_55 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09230_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\]
+ net855 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09161_ _04768_ _04769_ _04770_ _04771_ net786 net807 vssd1 vssd1 vccd1 vccd1 _04772_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__09254__A1 net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13050__A2 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ net756 _03623_ _03636_ _03638_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__and4_2
XFILLER_0_44_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09092_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1079 net1028 net1024 vssd1
+ vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__and4_2
XANTENNA__07937__B net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold900 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[964\] vssd1 vssd1
+ vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold911 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[452\] vssd1 vssd1
+ vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13889__B2 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[993\] vssd1 vssd1
+ vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\] vssd1 vssd1
+ vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[757\] vssd1 vssd1
+ vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[406\] vssd1 vssd1
+ vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\] vssd1 vssd1
+ vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[140\] vssd1 vssd1
+ vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_A _06073_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ net588 _05113_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__xnor2_1
Xhold988 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[151\] vssd1 vssd1
+ vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1017\] vssd1 vssd1
+ vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1118_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09644__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _04538_ _04544_ _04555_ net768 vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a22o_2
XANTENNA_fanout480_A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[48\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[16\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12864__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14786__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12077__B1 _07493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12616__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13813__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11824__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17341__1397 vssd1 vssd1 vccd1 vccd1 _17341__1397/HI net1397 sky130_fd_sc_hd__conb_1
X_09428_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[38\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[6\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09359_ _04966_ _04967_ _04968_ _04969_ net836 net749 vssd1 vssd1 vccd1 vccd1 _04970_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13041__A2 net382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ net236 net2608 net495 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__mux2_1
XANTENNA__08723__S net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11321_ net581 _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__or2_1
XANTENNA__10554__A team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_160_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14040_ net17 net1060 net1036 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] vssd1 vssd1
+ vccd1 vccd1 _01546_ sky130_fd_sc_hd__o22a_1
X_11252_ net553 _06663_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11369__B _06857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10203_ _03495_ net1055 _05809_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11937__X _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__A1 _07438_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11183_ _04166_ _04193_ net357 _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__o31a_1
XANTENNA__08959__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09554__S net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input41_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _05719_ _05744_ _05718_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ clknet_leaf_73_wb_clk_i _01667_ _00220_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15853__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13076__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10065_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] _04004_ vssd1
+ vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__nand2_1
X_14942_ net1239 vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__inv_2
XANTENNA__12855__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14873_ net1241 vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__inv_2
XANTENNA__14057__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16612_ clknet_leaf_171_wb_clk_i _02281_ _00841_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[585\]
+ sky130_fd_sc_hd__dfrtp_1
X_13824_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\] _05830_ net1099
+ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__mux2_1
XANTENNA__12607__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11815__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16543_ clknet_leaf_157_wb_clk_i _02212_ _00772_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[516\]
+ sky130_fd_sc_hd__dfrtp_1
X_13755_ _02992_ _03145_ _02994_ _02980_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__o211a_1
X_10967_ _04412_ _06291_ _06297_ net658 vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12706_ net2653 net407 net346 _07341_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a22o_1
X_16474_ clknet_leaf_39_wb_clk_i _02143_ _00703_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[447\]
+ sky130_fd_sc_hd__dfrtp_1
X_13686_ team_04_WB.MEM_SIZE_REG_REG\[0\] _03515_ net1046 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\]
+ _07685_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__o221a_1
X_10898_ net589 _06385_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13568__B1 _07697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15425_ net1130 vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12637_ _07608_ net488 net411 net2151 vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__a22o_1
XANTENNA__08039__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13032__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12568_ _07535_ net483 net417 net1708 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_152_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15356_ net1130 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Right_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ net2640 _03468_ _03470_ net818 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__o211a_1
X_11519_ _07007_ _07001_ _06997_ net465 vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_117_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12155__S net513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15287_ net1229 vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__inv_2
X_12499_ _07496_ net479 net424 net1829 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a22o_1
Xhold207 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\] vssd1 vssd1
+ vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[43\] vssd1 vssd1
+ vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\] vssd1 vssd1
+ vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ clknet_leaf_146_wb_clk_i _02695_ _01255_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_169_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14238_ _03426_ _03427_ net819 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_169_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12543__A1 net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13775__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[2\] _03385_
+ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and2_1
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13099__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08730_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[51\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[19\]
+ net870 vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__mux2_1
XANTENNA__12846__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1280 net1297 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_2
Xfanout1291 net1292 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__buf_4
X_08661_ _04266_ _04271_ net770 vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14048__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08592_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[52\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[20\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_52 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11267__D1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_191_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_165_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11461__C net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09213_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[10\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout326_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1068_A _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _04586_ _04644_ _04699_ _04754_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and4_1
XFILLER_0_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09075_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[620\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[588\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1235_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _03598_ _03609_ _03616_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__and3_2
Xhold730 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\] vssd1 vssd1
+ vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_536 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold741 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[581\] vssd1 vssd1
+ vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout695_A _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[449\] vssd1 vssd1
+ vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[450\] vssd1 vssd1
+ vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\] vssd1 vssd1
+ vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[541\] vssd1 vssd1
+ vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[736\] vssd1 vssd1
+ vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09374__S net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09227__X _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ net632 _04787_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout862_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[239\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[207\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_1
XANTENNA__12837__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout650_X net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ net731 _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or2_1
XANTENNA__14039__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11870_ _05466_ _07240_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10821_ _03808_ _06308_ net658 vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13540_ _02923_ _02929_ team_04_WB.ADDR_START_VAL_REG\[21\] vssd1 vssd1 vccd1 vccd1
+ _02931_ sky130_fd_sc_hd__a21oi_1
X_10752_ net573 _06207_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__or2_1
XANTENNA__09561__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__B1 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13471_ _02859_ _02861_ net997 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__mux2_1
X_10683_ team_04_WB.instance_to_wrap.final_design.uart.receiving _06159_ _06171_ vssd1
+ vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__and3_4
XFILLER_0_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09549__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15210_ net1107 vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__inv_2
X_12422_ net519 net601 _07386_ net432 net1734 vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a32o_1
XANTENNA__15140__A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16190_ clknet_leaf_157_wb_clk_i _01859_ _00419_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[163\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input89_A wbs_dat_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15848__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12773__A1 _07500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15141_ net1109 vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ net221 net670 vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__and2_2
XFILLER_0_106_875 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ _06546_ _06550_ net537 vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15072_ net1155 vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__inv_2
X_12284_ net229 net674 vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_75_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09077__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A1 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ _05338_ _05445_ _07235_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__or3_1
XANTENNA__13722__B1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_147_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ net571 _06647_ _06717_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_112_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ net706 _06651_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__o21a_1
XANTENNA__07952__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15959__CLK clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10117_ _05726_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__and2_1
X_15974_ clknet_leaf_51_wb_clk_i _01650_ _00203_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11097_ net635 net546 _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__a21bo_1
XANTENNA__12828__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10048_ _03591_ _04784_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nor2_1
X_14925_ net1152 vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_160_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[18\] vssd1 vssd1
+ vccd1 vccd1 net1527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11843__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ net1124 vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__inv_2
XANTENNA__08628__S net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ _03170_ _03195_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__o21a_1
XANTENNA__13789__B1 team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14787_ net1172 vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__inv_2
X_11999_ net219 net681 vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__and2_1
XANTENNA__11054__S net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16526_ clknet_leaf_27_wb_clk_i _02195_ _00755_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11264__A1 _04385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ net1001 _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or2_1
XANTENNA__12461__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16457_ clknet_leaf_120_wb_clk_i _02126_ _00686_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[430\]
+ sky130_fd_sc_hd__dfrtp_1
X_13669_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[0\] team_04_WB.MEM_SIZE_REG_REG\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_119_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13122__X _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15408_ net1173 vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16388_ clknet_leaf_167_wb_clk_i _02057_ _00617_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_756 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15339_ net1167 vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09900_ _03755_ _05508_ _05509_ _05510_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_20_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17009_ clknet_leaf_179_wb_clk_i _02678_ _01238_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09194__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout506 _07556_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__buf_4
X_17340__1396 vssd1 vssd1 vccd1 vccd1 _17340__1396/HI net1396 sky130_fd_sc_hd__conb_1
X_09831_ _03621_ _04611_ _04725_ _04784_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a31o_1
Xfanout517 _07449_ vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_6
Xfanout528 _06195_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_6
Xfanout539 net540 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
X_09762_ net732 _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or2_2
X_08713_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[755\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[723\]
+ net931 vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
X_09693_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[674\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\]
+ net888 vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__mux2_1
XANTENNA__13952__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08644_ net770 _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_174_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09791__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[630\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[598\]
+ net852 vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout443_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11255__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14128__X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout329_X net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09369__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_176_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_176_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_161_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09127_ _04734_ _04735_ _04736_ _04737_ net836 net748 vssd1 vssd1 vccd1 vccd1 _04738_
+ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1140_X net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10766__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09058_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[12\] team_04_WB.instance_to_wrap.CPU_DAT_O\[12\]
+ net1011 vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__mux2_4
XFILLER_0_130_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08009_ _03601_ _03603_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_92_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold560 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[83\] vssd1 vssd1
+ vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12523__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10832__A net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold571 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[611\] vssd1 vssd1
+ vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ team_04_WB.MEM_SIZE_REG_REG\[16\] _06508_ vssd1 vssd1 vccd1 vccd1 _06509_
+ sky130_fd_sc_hd__or2_1
Xhold582 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\] vssd1 vssd1
+ vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\] vssd1 vssd1
+ vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14023__B _05445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A1 net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10__f_wb_clk_i_A clknet_3_5_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07934__B2 _03535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__B net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ net610 _07341_ net474 net317 net1590 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a32o_1
XANTENNA__13207__X _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__A team_04_WB.MEM_SIZE_REG_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ net1224 vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__inv_2
X_11922_ net688 _07387_ _07388_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__a21oi_1
X_15690_ net1256 vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__inv_2
XANTENNA__12478__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14641_ net1267 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__inv_2
X_11853_ net757 _05878_ _06185_ _04387_ net689 vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10804_ net590 _04865_ _04919_ _04973_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__and4_1
X_14572_ net1286 vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__inv_2
X_11784_ net694 _07165_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16311_ clknet_leaf_166_wb_clk_i _01980_ _00540_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[284\]
+ sky130_fd_sc_hd__dfrtp_1
X_13523_ net1092 _02913_ net1043 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_64_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17291_ net1347 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10735_ _06220_ _06223_ net560 vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_902 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16242_ clknet_leaf_6_wb_clk_i _01911_ _00471_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[215\]
+ sky130_fd_sc_hd__dfrtp_1
X_13454_ team_04_WB.MEM_SIZE_REG_REG\[30\] _07871_ _02844_ vssd1 vssd1 vccd1 vccd1
+ _02845_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10666_ net1585 net1018 net1014 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1
+ vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ net1950 net432 _07630_ net519 vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
X_13385_ _07809_ _07810_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__nand2_1
X_16173_ clknet_leaf_43_wb_clk_i _01842_ _00402_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[146\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10597_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[1\]
+ _06136_ net1049 vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10221__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15124_ net1225 vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__clkbuf_4
X_12336_ net2231 net500 _07612_ net442 vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15055_ net1140 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__inv_2
X_12267_ net2440 net504 _07576_ net449 vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14006_ _05191_ _03336_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nor2_1
X_11218_ _06280_ _06703_ _06706_ net287 vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__o211a_1
X_12198_ net2508 net509 _07540_ net456 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_162_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09470__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__B1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _06272_ _06633_ _06635_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14120__B1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15957_ clknet_leaf_78_wb_clk_i _01633_ _00186_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13264__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12682__A0 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ net1128 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__inv_2
X_15888_ clknet_leaf_124_wb_clk_i _01565_ _00115_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__dfrtp_1
XANTENNA__08358__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14839_ net1229 vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__inv_2
XANTENNA__12956__X _07677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09978__A net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _03967_ _03968_ _03969_ _03970_ net828 net743 vssd1 vssd1 vccd1 vccd1 _03971_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16509_ clknet_leaf_131_wb_clk_i _02178_ _00738_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[482\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_160_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14095__S net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[187\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[155\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_926 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10917__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09189__S net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08093__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12691__X _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6__f_wb_clk_i_A clknet_3_3_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_20 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13947__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11960__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11748__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07945__B net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08169__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout303 _07681_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__buf_4
Xfanout314 _07677_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_4
Xfanout325 _07671_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout393_A _07672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_2
X_09814_ _05421_ _05422_ _05423_ _05424_ net834 net738 vssd1 vssd1 vccd1 vccd1 _05425_
+ sky130_fd_sc_hd__mux4_1
Xfanout347 net348 vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_4
Xfanout358 net359 vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1100_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[3\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout369 net372 vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14111__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\]
+ net902 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__mux2_1
XANTENNA__09669__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13465__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_905 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12673__A0 net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[162\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[130\]
+ net885 vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08627_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[564\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout825_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11770__X _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1188_X net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[502\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[470\]
+ net851 vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11779__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__A1 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ net770 _04093_ _04099_ net761 vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__A team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _06085_ net1544 net1020 vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10451_ _06025_ _06029_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__or2_1
XANTENNA__13925__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10203__A2 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13170_ _07606_ net382 net293 net2040 vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a22o_1
XANTENNA__11400__A1 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[6\] _05527_ vssd1
+ vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_131_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12121_ net2351 net354 _07515_ net455 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a22o_1
XANTENNA__11951__A2 _07075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12480__C net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ net2553 net517 _07479_ net455 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a22o_1
XANTENNA__09128__A net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 net133 vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08032__A _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _06317_ _06319_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_73_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_16860_ clknet_leaf_126_wb_clk_i _02529_ _01089_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[833\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09562__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_2
XANTENNA__14102__B1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout881 net882 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__buf_4
XANTENNA__15861__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_16791_ clknet_leaf_155_wb_clk_i _02460_ _01020_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout892 net894 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14309__A_N net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15742_ net1290 vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__inv_2
XANTENNA__12664__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12954_ net228 net2621 net320 vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__mux2_1
XANTENNA__09755__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\] vssd1 vssd1
+ vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14200__C net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ net652 net243 vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__and2_1
XFILLER_0_158_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15673_ net1258 vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _07585_ net345 net390 net1942 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22o_1
XANTENNA__12001__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output208_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11219__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ net1213 vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__inv_2
XANTENNA__10690__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ net2127 net526 net436 _07314_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a22o_1
XANTENNA__09507__S1 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12416__B1 net433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__S net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17343_ net1399 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14555_ net1179 vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11767_ net687 _07253_ _07254_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_155_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_155_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _02896_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__inv_2
X_17274_ net1333 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_10718_ net466 _05469_ _06201_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__or3_4
X_14486_ net1119 vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__inv_2
X_11698_ net585 _06946_ net288 vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16225_ clknet_leaf_133_wb_clk_i _01894_ _00454_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[198\]
+ sky130_fd_sc_hd__dfrtp_1
X_13437_ _07862_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__inv_2
X_10649_ _03542_ net1045 vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16156_ clknet_leaf_116_wb_clk_i _01825_ _00385_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[129\]
+ sky130_fd_sc_hd__dfrtp_1
X_13368_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08494__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13259__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ net1166 vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__inv_2
X_12319_ net260 net669 vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__and2_2
X_16087_ clknet_leaf_166_wb_clk_i _01756_ _00316_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_13299_ _06592_ net272 vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nand2_1
X_15038_ net1218 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09443__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14879__A net1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16989_ clknet_leaf_127_wb_clk_i _02658_ _01218_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12655__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ net588 net587 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and2_1
XANTENNA__08088__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09461_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[870\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[838\]
+ net888 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__mux2_1
X_08412_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[569\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[537\]
+ net843 vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__mux2_1
XANTENNA__10681__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09392_ net767 _05002_ _04991_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08816__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ _03950_ _03951_ _03952_ _03953_ net827 net744 vssd1 vssd1 vccd1 vccd1 _03954_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13080__A0 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09823__A1 _03634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10647__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_142 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08274_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[539\]
+ net929 vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout406_A _07664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13976__A_N _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09682__S0 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13686__A2 _03515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 net1110 vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_4
XANTENNA_fanout775_A net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12801__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12894__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__S net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout942_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] net1080 net1029 net1025 vssd1
+ vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11449__A1 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ net905 net754 _04782_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_87_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12646__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10672__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_191_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_191_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12670_ _07356_ net2484 net478 vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11621_ net565 _07063_ _07109_ net578 vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__o211ai_1
XANTENNA__13071__A0 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14029__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10557__A team_04_WB.instance_to_wrap.CPU_DAT_O\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ net1183 vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11621__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _05380_ net462 vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[1\] _03531_
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _06073_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14271_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[18\] _03447_
+ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__and2_1
X_11483_ net287 _06966_ _06971_ _06958_ net464 vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__a32o_2
XFILLER_0_52_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ clknet_leaf_52_wb_clk_i _01686_ _00239_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_150_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13222_ net79 team_04_WB.MEM_SIZE_REG_REG\[19\] net982 vssd1 vssd1 vccd1 vccd1 _01681_
+ sky130_fd_sc_hd__mux2_1
X_10434_ _06008_ _06010_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09557__S net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input71_A wbs_dat_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15856__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[10\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13079__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08250__A0 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ net279 _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__nor2_1
X_13153_ _07587_ net380 net296 net2166 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_5__f_wb_clk_i_X clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12104_ net251 net676 vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__and2_1
X_13084_ net232 net2424 net304 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__mux2_1
X_10296_ _05696_ _05756_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16912_ clknet_leaf_191_wb_clk_i _02581_ _01141_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\]
+ sky130_fd_sc_hd__dfrtp_1
X_12035_ net253 net680 vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12885__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09292__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11835__B net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16843_ clknet_leaf_16_wb_clk_i _02512_ _01072_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__B1 net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16774_ clknet_leaf_17_wb_clk_i _02443_ _01003_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13986_ _04641_ _03326_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_105_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12101__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15725_ net1295 vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12937_ _07333_ net2579 net319 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11851__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15656_ net1174 vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__inv_2
XANTENNA__10663__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _07568_ net332 net388 net2027 vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__a22o_1
X_14607_ net1282 vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__inv_2
XANTENNA__13062__A0 _07283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11819_ net704 _05832_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_174_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08608__A2 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15587_ net1170 vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12158__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_174_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12799_ net239 net2586 net322 vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17326_ net1382 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ net1285 vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_79 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17257_ net1317 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XANTENNA__13778__A team_04_WB.ADDR_START_VAL_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09018__C1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14469_ net1250 vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16208_ clknet_leaf_3_wb_clk_i _01877_ _00437_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[181\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09467__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12168__A2 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17188_ clknet_leaf_87_wb_clk_i _02800_ _01417_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ clknet_leaf_23_wb_clk_i _01808_ _00368_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13117__A1 _07549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09991__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\]
+ net880 vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_1
XANTENNA__09416__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07912_ net1101 net1080 vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nand2_1
XANTENNA__12876__B1 net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08892_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[368\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[336\]
+ net873 vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__mux2_1
XANTENNA__10930__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__C net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12628__B1 net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09513_ _05120_ _05121_ _05122_ _05123_ net832 net737 vssd1 vssd1 vccd1 vccd1 _05124_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13960__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__A0 _05475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1098_A team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15233__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__A2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ _05049_ _05054_ net775 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__mux2_1
XANTENNA__08546__S net918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1071 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_166_Right_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09375_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[167\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[135\]
+ net945 vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__mux2_1
XANTENNA__13053__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1265_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08155__S0 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12800__A0 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08326_ _03933_ _03934_ _03935_ _03936_ net788 net809 vssd1 vssd1 vccd1 vccd1 _03937_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11603__A1 _05219_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08257_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[315\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09377__S net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08188_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[540\]
+ net876 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout892_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A2 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1220_X net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_103_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _05690_ _05691_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[18\] _04387_ vssd1
+ vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12531__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786__5 clknet_leaf_75_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08630__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _03228_ _03230_ _02855_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__a21o_1
XANTENNA__12619__B1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13771_ _07829_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__and2_1
X_10983_ _06466_ _06471_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__and2_1
XANTENNA__12095__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15510_ net1223 vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ net2172 net406 net345 _07439_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16490_ clknet_leaf_164_wb_clk_i _02159_ _00719_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ net1274 vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13044__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ _06191_ _06194_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__or2_4
XFILLER_0_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ _05219_ net578 net358 _07092_ net462 vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__o311a_1
XFILLER_0_26_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15372_ net1129 vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_142_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12584_ _07551_ net490 net418 net2033 vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a22o_1
X_17111_ clknet_leaf_104_wb_clk_i _02746_ _01340_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08697__S1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[15\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[14\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[13\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[12\] net1091
+ net1089 vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__mux4_1
XFILLER_0_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11535_ net754 _07023_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__and2_1
XANTENNA__08471__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17042_ clknet_leaf_9_wb_clk_i _02711_ _01271_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
X_14254_ _03437_ net819 _03436_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__and3b_1
X_11466_ net753 _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__nand2_2
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09646__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ _03518_ net1072 _07699_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_78_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10417_ net1090 net1089 _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_78_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14185_ _03373_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11397_ _05464_ _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__nor2_2
XANTENNA__12007__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08774__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ _07570_ net373 net295 net1890 vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__a22o_1
XANTENNA__12570__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10348_ net623 _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__nor2_1
X_10279_ _05639_ net622 _05873_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a31o_1
X_13067_ net237 net2549 net302 vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__mux2_1
XANTENNA__12858__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12322__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ net2593 net516 _07462_ net448 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11530__B1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16826_ clknet_leaf_44_wb_clk_i _02495_ _01055_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16757_ clknet_leaf_31_wb_clk_i _02426_ _00986_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09487__C1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ net1668 net1069 _03318_ net264 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_181_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13272__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ net1281 vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__inv_2
XANTENNA__11833__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16688_ clknet_leaf_191_wb_clk_i _02357_ _00917_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[661\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12396__B net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10909__B _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15639_ net1177 vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_67 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13035__B1 net306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13586__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[939\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[907\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13586__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09254__A2 _04864_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ net759 _03622_ _03635_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__or3_1
X_17309_ net1365 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09197__S net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1078 net1030 net1026 vssd1
+ vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_77 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_99 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold901 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[772\] vssd1 vssd1
+ vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\] vssd1 vssd1
+ vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold923 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[466\] vssd1 vssd1
+ vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[810\] vssd1 vssd1
+ vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[536\] vssd1 vssd1
+ vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[847\] vssd1 vssd1
+ vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__A2 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold967 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[908\] vssd1 vssd1
+ vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[415\] vssd1 vssd1
+ vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ net588 _05113_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__and2b_1
Xhold989 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[945\] vssd1 vssd1
+ vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ _04549_ _04554_ net774 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__mux2_1
XANTENNA__12849__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[80\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09660__S net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__A0 net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12077__B2 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09427_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[102\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[70\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13026__B1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout526_X net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08128__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__A _03781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09358_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[936\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[904\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08309_ _03892_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09289_ net721 _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__or2_1
XANTENNA__12526__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ net575 _06534_ _06807_ _06804_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__o31a_1
XFILLER_0_105_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ net535 _06527_ _06528_ net558 vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_160_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ net277 _05808_ _05807_ net1074 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ net592 _04193_ net360 vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10133_ _05722_ _05743_ _05721_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_73_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15138__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ clknet_leaf_79_wb_clk_i _01666_ _00219_ vssd1 vssd1 vccd1 vccd1 team_04_WB.MEM_SIZE_REG_REG\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_73_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13501__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12304__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13501__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[25\] _04004_ vssd1
+ vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__or2_1
XANTENNA_input34_A gpio_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ net1155 vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__inv_2
X_14872_ net1205 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__inv_2
XANTENNA__08975__A _04557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16611_ clknet_leaf_125_wb_clk_i _02280_ _00840_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[584\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13265__A0 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13823_ net1092 _03213_ net1043 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[24\]
+ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_49 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17309__1365 vssd1 vssd1 vccd1 vccd1 _17309__1365/HI net1365 sky130_fd_sc_hd__conb_1
X_16542_ clknet_leaf_142_wb_clk_i _02211_ _00771_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[515\]
+ sky130_fd_sc_hd__dfrtp_1
X_13754_ _03109_ _03119_ _03122_ _03144_ _03108_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o221a_1
XANTENNA__08186__S net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10966_ _06291_ _06297_ net658 vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12705_ net2045 net405 net335 _07334_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a22o_1
X_16473_ clknet_leaf_178_wb_clk_i _02142_ _00702_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[446\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13017__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ team_04_WB.MEM_SIZE_REG_REG\[0\] net993 net991 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\]
+ net1000 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__o221a_1
X_10897_ _05003_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15424_ net1212 vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12636_ _07607_ net484 net409 net1653 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08914__S net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__A3 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15355_ net1112 vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__inv_2
XFILLER_0_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12567_ _07534_ net484 net417 net1891 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10745__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\] _03468_
+ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11518_ _06833_ _07006_ net583 vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15286_ net1221 vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_117_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12498_ _07495_ net479 net424 net1718 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold208 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\] vssd1 vssd1
+ vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17025_ clknet_leaf_133_wb_clk_i _02694_ _01254_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold219 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[574\] vssd1 vssd1
+ vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14237_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[3\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ _03422_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\] vssd1 vssd1
+ vccd1 vccd1 _03427_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_148 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11449_ _04557_ net635 net546 vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_169_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_169_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09745__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ _03385_ _03386_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[1\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08502__X _04113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__S net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ _07551_ net378 net300 net1856 vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_84_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14099_ net1 _07701_ _07699_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a21o_1
XANTENNA__09172__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout1270 net1279 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__buf_4
Xfanout1281 net1288 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__buf_4
X_08660_ _04267_ _04268_ _04269_ _04270_ net783 net805 vssd1 vssd1 vccd1 vccd1 _04271_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_1_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1292 net1293 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__buf_4
XFILLER_0_89_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13256__A0 net81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16809_ clknet_leaf_99_wb_clk_i _02478_ _01038_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[782\]
+ sky130_fd_sc_hd__dfrtp_1
X_08591_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[116\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[84\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11806__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_751 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13008__B1 net312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09212_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[106\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[74\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08824__S net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09143_ _04724_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12231__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11103__X _06592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_A _07675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12782__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ _03597_ _03607_ _03617_ _03625_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold720 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[471\] vssd1 vssd1
+ vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[803\] vssd1 vssd1
+ vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[293\] vssd1 vssd1
+ vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09655__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold753 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\] vssd1 vssd1
+ vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11757__Y _07246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold764 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[175\] vssd1 vssd1
+ vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[222\] vssd1 vssd1
+ vccd1 vccd1 net2212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[998\] vssd1 vssd1
+ vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\] vssd1 vssd1
+ vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ net634 _04671_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ net776 _04537_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or2_1
XANTENNA__12298__B2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08858_ _04465_ _04466_ _04467_ _04468_ net837 net748 vssd1 vssd1 vccd1 vccd1 _04469_
+ sky130_fd_sc_hd__mux4_1
X_08789_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[882\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[850\]
+ net869 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ net658 _06308_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__or2_1
XANTENNA__12110__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15802__21 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12470__A1 net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10751_ net577 _06207_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_98_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13470_ net994 _02858_ _02860_ net989 vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clknet_4_6__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10682_ _06159_ _06171_ _03517_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_164_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13014__A3 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12421_ net521 net605 _07381_ net433 net1631 vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a32o_1
XFILLER_0_152_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12222__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12773__A2 net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ net1188 vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__inv_2
X_12352_ net2168 net501 _07620_ net456 vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__B1 net457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11303_ _06791_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15071_ net1270 vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__inv_2
X_12283_ net2383 net505 _07584_ net451 vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09077__S1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022_ _07688_ net1041 _03347_ net1072 net1491 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__a32o_1
XANTENNA__09418__X _05029_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__S net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11234_ net289 _06719_ _06720_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15864__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_X clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13087__S net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] _05113_ vssd1
+ vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__or2_1
X_15973_ clknet_leaf_50_wb_clk_i _01649_ _00202_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_11096_ _04724_ net552 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__nand2_1
XANTENNA__12289__B2 net455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ net646 _03646_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08588__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14924_ net1121 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__inv_2
XANTENNA__11497__C1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 net109 vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_160_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_160_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 net141 vssd1 vssd1 vccd1 vccd1 net1528 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13238__A0 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__B net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14855_ net1142 vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__inv_2
X_13806_ _03157_ _03196_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__C net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14786_ net1255 vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__inv_2
X_11998_ net2305 net517 _07452_ net450 vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
X_16525_ clknet_leaf_40_wb_clk_i _02194_ _00754_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[498\]
+ sky130_fd_sc_hd__dfrtp_1
X_13737_ net995 _03124_ _03127_ net991 vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10949_ _05462_ _06287_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__nand2_1
XANTENNA__12461__A1 net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16456_ clknet_leaf_113_wb_clk_i _02125_ _00685_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\]
+ sky130_fd_sc_hd__dfrtp_1
X_13668_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[2\] net1102 vssd1
+ vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_119_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13005__A3 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14202__A2 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ net1195 vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__inv_2
X_12619_ _07588_ net493 net415 net2053 vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22o_1
X_16387_ clknet_leaf_121_wb_clk_i _02056_ _00616_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[360\]
+ sky130_fd_sc_hd__dfrtp_1
X_13599_ team_04_WB.ADDR_START_VAL_REG\[12\] _02989_ vssd1 vssd1 vccd1 vccd1 _02990_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10224__B1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15338_ net1112 vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__inv_2
XANTENNA__12764__A2 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13961__A1 _03973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15269_ net1108 vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__inv_2
XANTENNA__12690__A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17008_ clknet_leaf_192_wb_clk_i _02677_ _01237_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[981\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12516__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09830_ _04611_ _04725_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_8
Xfanout518 _07449_ vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_2
Xfanout529 _06195_ vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__buf_2
X_09761_ _05368_ _05369_ _05370_ _05371_ net837 net749 vssd1 vssd1 vccd1 vccd1 _05372_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__08111__C _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__X _07082_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08712_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[563\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[531\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__mux2_1
X_09692_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[738\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[706\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__mux2_1
XANTENNA__08819__S net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13229__A0 net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _04250_ _04251_ _04252_ _04253_ net783 net800 vssd1 vssd1 vccd1 vccd1 _04254_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08574_ _04181_ _04182_ _04183_ _04184_ net825 net742 vssd1 vssd1 vccd1 vccd1 _04185_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10369__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_423 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout436_A net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08554__S net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12204__B2 net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout603_A net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12755__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[429\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[397\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10766__A1 net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ net765 _04667_ _04656_ _04655_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_170_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12804__S net323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ _03601_ _03603_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__a211oi_1
XANTENNA__12507__A2 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17308__1364 vssd1 vssd1 vccd1 vccd1 _17308__1364/HI net1364 sky130_fd_sc_hd__conb_1
XFILLER_0_163_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_145_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold550 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[616\] vssd1 vssd1
+ vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[680\] vssd1 vssd1
+ vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_A _03555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold572 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\] vssd1 vssd1
+ vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[889\] vssd1 vssd1
+ vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13180__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[619\] vssd1 vssd1
+ vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10551__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__B1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _04329_ _04331_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ net604 _07334_ net470 net315 net1586 vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a32o_1
XANTENNA__12140__A0 _07333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11921_ _03631_ _05947_ _05949_ net760 net695 vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__a221o_1
XANTENNA__11494__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12478__C net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14640_ net1175 vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11852_ net2300 net527 net447 _07328_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ net659 _06286_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14571_ net1286 vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11783_ _03631_ _05795_ net694 _07268_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_1038 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12443__B2 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16310_ clknet_leaf_10_wb_clk_i _01979_ _00539_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[283\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_99_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13522_ _07846_ _02912_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__or2_1
XANTENNA__08742__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17290_ net1346 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XANTENNA__12994__A2 net470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10734_ _06221_ _06222_ net538 vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__mux2_1
XANTENNA__08464__S net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15859__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ clknet_leaf_172_wb_clk_i _01910_ _00470_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\]
+ sky130_fd_sc_hd__dfrtp_1
X_13453_ _07871_ _02842_ _02843_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__nor3_1
XFILLER_0_125_426 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ net1518 net1018 net1014 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1
+ vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_149_Left_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12404_ net651 net600 net241 vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__and3_1
XANTENNA__12746__A2 net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16172_ clknet_leaf_107_wb_clk_i _01841_ _00401_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[145\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13384_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] team_04_WB.MEM_SIZE_REG_REG\[9\]
+ _07808_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__or3_1
XANTENNA__09072__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] net1096 net1051 vssd1 vssd1 vccd1
+ vccd1 _06136_ sky130_fd_sc_hd__and3_1
XFILLER_0_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09611__A2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15123_ net1233 vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12335_ net254 net669 vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__and2_2
XFILLER_0_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15054_ net1197 vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__inv_2
X_12266_ net243 net672 vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14005_ _05083_ net265 _03335_ _03338_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13171__A2 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ net640 _04030_ net357 _06704_ _06705_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__o311a_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12015__A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ net255 net650 vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__and2_1
XANTENNA__11182__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_162_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09470__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11148_ net572 _06636_ net581 vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21o_1
XANTENNA__13459__B1 _02846_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_158_Left_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14120__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__B2 team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15956_ clknet_leaf_79_wb_clk_i _01632_ _00185_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11079_ net625 net547 vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__nand2_1
X_14907_ net1126 vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__inv_2
X_15887_ clknet_leaf_123_wb_clk_i _01564_ _00114_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11890__C1 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14838_ net1222 vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14769_ net1265 vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15061__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793__12 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__inv_2
XANTENNA__12985__A2 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16508_ clknet_leaf_128_wb_clk_i _02177_ _00737_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08374__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[251\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[219\]
+ net863 vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_167_Left_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_938 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ clknet_leaf_167_wb_clk_i _02108_ _00668_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[412\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09994__A net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12737__A2 net336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10748__A1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13162__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 net305 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12370__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__A1 _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout315 _07677_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_4
Xfanout326 net332 vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_4
Xfanout337 _07667_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_2
X_09813_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\]
+ net893 vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__mux2_1
Xfanout348 net349 vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_2
XANTENNA__10920__A1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 _06258_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout386_A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ net748 _05354_ net726 vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09675_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[226\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10684__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[628\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[596\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10099__B _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _04167_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__inv_2
XANTENNA__12425__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout720_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08284__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ net779 _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__or2_1
XANTENNA__10987__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_730 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12728__A2 net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10450_ _06023_ _06027_ _06024_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09109_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[685\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[653\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__mux2_1
XANTENNA__08801__A0 _04387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _05722_ _05743_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_131_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12534__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12120_ net228 net678 vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__and2_1
XFILLER_0_130_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12051_ net221 net683 vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__and2_1
XANTENNA__13153__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[417\] vssd1 vssd1
+ vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\] vssd1 vssd1
+ vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08032__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _06324_ _06489_ _06319_ _06322_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12900__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
Xfanout871 net904 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__buf_2
Xfanout882 net883 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__clkbuf_4
X_16790_ clknet_leaf_15_wb_clk_i _02459_ _01019_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_4
X_15741_ net1284 vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__inv_2
X_12953_ net221 net2606 net321 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__mux2_1
XANTENNA__13861__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1080 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\] vssd1 vssd1
+ vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1091 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[519\] vssd1 vssd1
+ vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ net694 _06972_ _07373_ net615 vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_107_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15672_ net1262 vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_42_wb_clk_i clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_66_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _07584_ net341 net390 net1934 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a22o_1
X_14623_ net1241 vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ net651 net236 vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__and2_1
XANTENNA__12416__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output103_A net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17342_ net1398 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XANTENNA__08715__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14554_ net1179 vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__inv_2
XANTENNA__12967__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11766_ net757 _05784_ _06185_ _03728_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10737__B net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ team_04_WB.ADDR_START_VAL_REG\[26\] _02894_ vssd1 vssd1 vccd1 vccd1 _02896_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_155_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17273_ net1332 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10717_ _05473_ net465 vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__or2_2
X_14485_ net1163 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11697_ _06331_ _06487_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ clknet_leaf_140_wb_clk_i _01893_ _00453_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[197\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12719__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13436_ _07860_ _07861_ _07728_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__o21a_1
X_10648_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\] net1081
+ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__nand2_1
XANTENNA__08922__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09596__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11849__A net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16155_ clknet_leaf_104_wb_clk_i _01824_ _00384_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[128\]
+ sky130_fd_sc_hd__dfrtp_1
X_13367_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] team_04_WB.MEM_SIZE_REG_REG\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_98_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10579_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[7\]
+ _06124_ net1049 vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15106_ net1265 vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__inv_2
X_12318_ net2124 net499 _07603_ net437 vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a22o_1
X_16086_ clknet_leaf_18_wb_clk_i _01755_ _00315_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_13298_ _07719_ _07718_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13144__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15037_ net1154 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__inv_2
X_12249_ net2384 net503 _07567_ net436 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11155__A1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__S net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__B1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13275__S net978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16988_ clknet_leaf_127_wb_clk_i _02657_ _01217_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[961\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_147_Right_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15939_ clknet_leaf_52_wb_clk_i _01616_ _00166_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dfrtp_1
XANTENNA__14895__A net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11871__X _07345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10666__B1 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ net731 _05070_ net714 vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__o21a_1
XFILLER_0_171_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08411_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[633\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[601\]
+ net844 vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09391_ _04996_ _05001_ net774 vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__mux2_1
XANTENNA__12407__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17307__1363 vssd1 vssd1 vccd1 vccd1 _17307__1363/HI net1363 sky130_fd_sc_hd__conb_1
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12958__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08342_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[186\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[154\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10647__B _06174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09823__A2 _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08273_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[635\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[603\]
+ net929 vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13958__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout301_A _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1043_A net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12591__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__S1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09229__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13135__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1210_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout670_A _07589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_X net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout389_X net389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07988_ _03512_ _03547_ _03593_ _03595_ _03596_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09727_ net905 net754 vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nand2_1
XANTENNA__09198__S0 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout935_A net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12102__B net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__B1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _05265_ _05266_ _05267_ _05268_ net794 net803 vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_26_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[500\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[468\]
+ net842 vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12529__S net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ _05196_ _05197_ _05198_ _05199_ net794 net814 vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10838__A _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ net533 _07096_ _07108_ net556 vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14029__B team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_132_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _07025_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ net2635 _06000_ _06051_ _03521_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
X_14270_ _03447_ net820 _03446_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__and3b_1
XANTENNA__14020__B1 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11482_ _04699_ net365 _06969_ _06970_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__o211a_1
XFILLER_0_107_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_160_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_160_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_162_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13674__A1_N net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11909__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ net81 team_04_WB.MEM_SIZE_REG_REG\[20\] net982 vssd1 vssd1 vccd1 vccd1 _01682_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09122__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10433_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[8\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\]
+ _03528_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_150_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12582__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__B2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input64_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _07586_ net378 net297 net2042 vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__a22o_1
X_10364_ _05529_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__nor2_1
XANTENNA__08250__A1 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08043__A team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12103_ net2061 net352 _07506_ net442 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13126__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ net223 net2524 net304 vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__mux2_1
X_10295_ _05577_ _05636_ net624 _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__o211a_1
XANTENNA__12334__B1 _07611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16911_ clknet_leaf_188_wb_clk_i _02580_ _01140_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[884\]
+ sky130_fd_sc_hd__dfrtp_1
X_12034_ net2400 net515 _07470_ net442 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a22o_1
XANTENNA__15872__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[26\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_109_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16842_ clknet_leaf_160_wb_clk_i _02511_ _01071_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09750__B2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout690 net692 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__buf_2
XFILLER_0_137_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16773_ clknet_leaf_4_wb_clk_i _02442_ _01002_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[746\]
+ sky130_fd_sc_hd__dfrtp_1
X_13985_ net1572 net1070 _03327_ net265 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_171_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_15724_ net1294 vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__inv_2
XANTENNA__11845__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ net2613 net319 _07676_ net260 vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__a22o_1
XANTENNA__15604__A net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ net1174 vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _07567_ net326 net388 net2093 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14606_ net1281 vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__inv_2
X_11818_ net686 _07298_ _07297_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15586_ net1219 vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ net241 net2372 net322 vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ net1381 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
X_14537_ net1263 vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__inv_2
X_11749_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[7\]
+ net274 vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09748__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17256_ net1316 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XFILLER_0_148_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08652__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14468_ net1250 vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_896 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13419_ _07745_ _07840_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__a21oi_1
X_16207_ clknet_leaf_186_wb_clk_i _01876_ _00436_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\]
+ sky130_fd_sc_hd__dfrtp_1
X_17187_ clknet_leaf_88_wb_clk_i _02799_ _01416_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_14399_ net1283 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12573__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16138_ clknet_leaf_109_wb_clk_i _01807_ _00367_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13117__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16069_ clknet_leaf_6_wb_clk_i _01738_ _00298_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_08960_ net731 _04564_ net715 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09416__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09483__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ team_04_WB.instance_to_wrap.BUSY_O net1101 team_04_WB.EN_VAL_REG vssd1 vssd1
+ vccd1 vccd1 _03525_ sky130_fd_sc_hd__and3b_1
XANTENNA__09336__X _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ _03558_ net702 _04386_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a21oi_2
XANTENNA__08099__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07942__D net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12203__A net253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[36\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[4\]
+ net879 vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__mux2_1
XANTENNA__07911__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _05050_ _05051_ _05052_ _05053_ net793 net802 vssd1 vssd1 vccd1 vccd1 _05054_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout251_A net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout349_A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09374_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[231\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[199\]
+ net952 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08155__S1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[954\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[922\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout516_A _07449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1258_A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10811__B1 net658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08256_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[379\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[347\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08187_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[636\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[604\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12564__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout885_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13108__A2 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12812__S net322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\] _04331_ vssd1
+ vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_89_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08091__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_113_Left_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11952__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15424__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13770_ _07750_ _07825_ _07828_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__or3b_1
XANTENNA__11827__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _04501_ _06356_ _06465_ _04440_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12095__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12721_ net2156 net406 net344 _07433_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15440_ net1164 vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _07623_ net493 net411 net1774 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13044__A1 _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11603_ _05219_ net578 net361 vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__a21o_1
X_15371_ net1167 vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_152_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _07550_ net489 net418 net2008 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14322_ net1087 _03478_ _03481_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a211o_1
X_17110_ clknet_leaf_91_wb_clk_i _02745_ _01339_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07877__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11534_ net462 _07012_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15867__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[21\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Left_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17041_ clknet_leaf_179_wb_clk_i _02710_ _01270_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14253_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ _03433_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__and3_1
XFILLER_0_162_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10507__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11465_ _06206_ _06945_ _06953_ _06936_ net462 vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__o32a_2
X_13204_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__or2_1
XANTENNA__12555__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__S1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[0\] net1088
+ net1087 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__and4b_1
XFILLER_0_111_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\]
+ _03393_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08223__B2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11396_ net583 _06250_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__nand2_2
XFILLER_0_150_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ _07569_ net373 net295 net1997 vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a22o_1
X_10347_ _05713_ _05749_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17306__1362 vssd1 vssd1 vccd1 vccd1 _17306__1362/HI net1362 sky130_fd_sc_hd__conb_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13066_ net248 net2243 net303 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__mux2_1
X_10278_ net622 _05875_ net277 vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__o21ai_1
X_12017_ net260 net681 vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__and2_1
XANTENNA__10869__B1 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12023__A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16825_ clknet_leaf_151_wb_clk_i _02494_ _01054_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[798\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_124_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16756_ clknet_leaf_3_wb_clk_i _02425_ _00985_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[729\]
+ sky130_fd_sc_hd__dfrtp_1
X_13968_ _04192_ net599 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__and2b_2
X_15707_ net1281 vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12919_ _07621_ net344 net387 net1777 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a22o_1
X_13899_ _03182_ _03190_ _03274_ net1042 vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__o31a_1
X_16687_ clknet_leaf_189_wb_clk_i _02356_ _00916_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12396__C net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15638_ net1178 vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09334__S0 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15569_ net1271 vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__inv_2
XANTENNA__12794__A0 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08110_ net766 _03720_ _03709_ _03703_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09478__S net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17308_ net1364 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
XFILLER_0_173_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09090_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\]
+ net965 vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08041_ team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] net1079 net1028 net1024 vssd1
+ vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__and4b_2
X_17239_ net1300 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_25_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold902 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[740\] vssd1 vssd1
+ vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11102__A _05473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold913 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[990\] vssd1 vssd1
+ vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A2 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold924 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\] vssd1 vssd1
+ vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\] vssd1 vssd1
+ vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[836\] vssd1 vssd1
+ vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold957 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\] vssd1 vssd1
+ vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\] vssd1 vssd1
+ vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09992_ _05601_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__and2_1
Xhold979 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[933\] vssd1 vssd1
+ vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap698 _05453_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08943_ _04550_ _04551_ _04552_ _04553_ net792 net812 vssd1 vssd1 vccd1 vccd1 _04554_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout299_A _07682_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13510__A2 net272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[176\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11809__C1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12077__A2 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08376__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09573__S0 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10388__A net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout633_A _04779_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ _05033_ _05034_ _05035_ _05036_ net793 net813 vssd1 vssd1 vccd1 vccd1 _05037_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08128__S1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09357_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[968\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12807__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09388__S net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12785__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08308_ _03894_ _03918_ net663 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__mux2_2
XANTENNA__08292__S net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_362 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09288_ _04895_ _04896_ _04897_ _04898_ net826 net734 vssd1 vssd1 vccd1 vccd1 _04899_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08239_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[829\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__A _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10554__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ net553 _06736_ _06737_ _06735_ net572 vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__o311a_1
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10201_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _05541_ vssd1
+ vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08300__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _06669_ _06668_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10851__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10132_ _05724_ _05742_ _05723_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10063_ _05672_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__nor2_1
X_14940_ net1127 vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A DAT_I[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ net1226 vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__inv_2
X_16610_ clknet_leaf_149_wb_clk_i _02279_ _00839_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11682__A net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13822_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13753_ _03131_ _03140_ _03130_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a21oi_1
X_16541_ clknet_leaf_132_wb_clk_i _02210_ _00770_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10965_ _06445_ _06453_ _06357_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11815__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ net1831 net405 net336 _07328_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ net274 _07058_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__and2b_1
X_16472_ clknet_leaf_151_wb_clk_i _02141_ _00701_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[445\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ _05030_ _06384_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xor2_1
XANTENNA__13568__A2 net273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12635_ _07606_ net493 net410 net1743 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a22o_1
X_15423_ net1273 vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Left_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12776__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15354_ net1146 vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08444__A1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ _07533_ net479 net416 net2140 vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14305_ _03468_ _03469_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ net577 _07004_ _07005_ _06251_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ net1209 vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__inv_2
X_12497_ _07494_ net481 net424 net1806 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14236_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[5\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\]
+ _03423_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17024_ clknet_leaf_135_wb_clk_i _02693_ _01253_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[997\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold209 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[695\] vssd1 vssd1
+ vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ _06247_ _06746_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08930__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11200__A0 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_169_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14167_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\] _03383_
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__o21ai_1
X_11379_ _06364_ _06866_ net464 vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__o21a_1
X_13118_ _07550_ net379 net300 net1858 vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__a22o_1
X_14098_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\] _07688_ _07694_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\]
+ _03516_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a32o_1
XANTENNA__08231__A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ _07510_ net378 net308 net1621 vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__a22o_1
Xfanout1260 net1261 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12700__B1 net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1271 net1279 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__buf_2
Xfanout1282 net1288 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12688__A net614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1293 net1297 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__clkbuf_2
X_16808_ clknet_leaf_114_wb_clk_i _02477_ _01037_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[781\]
+ sky130_fd_sc_hd__dfrtp_1
X_08590_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[180\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[148\]
+ net909 vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16739_ clknet_leaf_122_wb_clk_i _02408_ _00968_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11806__A2 _06708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10001__A _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13008__A1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[170\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[138\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12767__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09142_ _04727_ _04752_ net666 vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__mux2_2
XANTENNA__12231__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09073_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\]
+ net854 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout214_A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12519__B1 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _03625_ _03608_ _03598_ _03616_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__and4b_4
XFILLER_0_13_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold710 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[819\] vssd1 vssd1
+ vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13966__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold721 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[348\] vssd1 vssd1
+ vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\] vssd1 vssd1
+ vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold743 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[946\] vssd1 vssd1
+ vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12362__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12215__X _07549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold754 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[763\] vssd1 vssd1
+ vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[823\] vssd1 vssd1
+ vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08294__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1123_A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[580\] vssd1 vssd1
+ vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[566\] vssd1 vssd1
+ vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _04723_ _04728_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__or2_1
Xhold798 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[691\] vssd1 vssd1
+ vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ _04533_ _04534_ _04535_ _04536_ net798 net817 vssd1 vssd1 vccd1 vccd1 _04537_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13982__A _07344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12298__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[689\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15970__Q team_04_WB.ADDR_START_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_X net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13247__A1 team_04_WB.ADDR_START_VAL_REG\[29\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ net729 _04392_ net713 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08287__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1280_X net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout636_X net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15702__A net1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10750_ _06233_ _06238_ net560 vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12470__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[999\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__mux2_1
XANTENNA__09700__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17305__1361 vssd1 vssd1 vccd1 vccd1 _17305__1361/HI net1361 sky130_fd_sc_hd__conb_1
XFILLER_0_138_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10681_ net1628 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1
+ vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12537__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12758__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ net522 net606 _07375_ net432 net1709 vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a32o_1
XFILLER_0_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08390__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12222__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_164_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12351_ net230 net670 vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__and2_2
XFILLER_0_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_67_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _06543_ _06586_ net531 vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__mux2_1
X_15070_ net1218 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__inv_2
X_12282_ net231 net674 vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ _07345_ _03345_ _07694_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__a21o_1
XANTENNA__13183__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ net585 _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__nand2_1
XANTENNA__10581__A team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12930__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ _06516_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_112_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14132__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_164_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10115_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] _05113_ vssd1
+ vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_164_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15972_ clknet_leaf_50_wb_clk_i _01648_ _00201_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12289__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ net632 net552 _06583_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__a21bo_1
XANTENNA__08986__A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ _05548_ _05655_ _05546_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__a21o_1
XANTENNA__08588__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14923_ net1162 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_160_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[28\]
+ vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[16\] vssd1 vssd1
+ vccd1 vccd1 net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 net125 vssd1 vssd1 vccd1 vccd1 net1529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10520__S net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08197__S net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14854_ net1108 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__inv_2
X_13805_ team_04_WB.ADDR_START_VAL_REG\[19\] _03156_ _03168_ vssd1 vssd1 vccd1 vccd1
+ _03196_ sky130_fd_sc_hd__o21a_1
X_11997_ net214 net682 vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__and2_1
X_14785_ net1150 vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__inv_2
XANTENNA__08114__B1 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12997__B1 net310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ clknet_leaf_112_wb_clk_i _02193_ _00753_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[497\]
+ sky130_fd_sc_hd__dfrtp_1
X_13736_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05949_ net1102
+ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
X_10948_ _06432_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nor2_1
XANTENNA__08925__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__A2 net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__A3 _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16455_ clknet_leaf_24_wb_clk_i _02124_ _00684_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\]
+ sky130_fd_sc_hd__dfrtp_1
X_13667_ net274 _07693_ _07090_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__or3b_1
X_10879_ _06362_ _06363_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__or3b_1
XFILLER_0_112_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12749__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15406_ net1203 vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12618_ _07587_ net491 net414 net2519 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13598_ net999 _02985_ _02988_ _02983_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16386_ clknet_leaf_146_wb_clk_i _02055_ _00615_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[359\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08417__B2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11421__A0 net635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15337_ net1137 vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__inv_2
X_12549_ net2106 net231 net422 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
XANTENNA__13961__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11972__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15268_ net1188 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__inv_2
XFILLER_0_123_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10762__Y _06251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13174__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11587__A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17007_ clknet_leaf_189_wb_clk_i _02676_ _01236_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\]
+ sky130_fd_sc_hd__dfrtp_1
X_14219_ _06051_ _06074_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.next_state\[0\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_112_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15199_ net1250 vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__inv_2
XANTENNA__12921__B1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 net510 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_8
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_4
X_09760_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[672\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\]
+ net901 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__mux2_1
XANTENNA__13477__B2 net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[627\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[595\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__mux2_1
XANTENNA__08579__S1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[546\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[514\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__mux2_1
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
X_08642_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[309\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[277\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__mux2_1
XANTENNA__12211__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[950\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[918\]
+ net851 vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__B1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13684__A_N net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout331_A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_A _07700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout429_A _07641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12204__A2 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09125_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[493\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[461\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11963__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09056_ _04661_ _04666_ net773 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08570__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ _03598_ _03616_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nand2_1
XANTENNA__13165__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout798_A net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold540 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[874\] vssd1 vssd1
+ vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold551 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[545\] vssd1 vssd1
+ vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12912__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\] vssd1 vssd1
+ vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[221\] vssd1 vssd1
+ vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold584 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[364\] vssd1 vssd1
+ vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\] vssd1 vssd1
+ vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout965_A net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14114__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__S net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_185_wb_clk_i clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_185_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_142_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[624\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[592\]
+ net864 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _04385_ _04412_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_114_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_11920_ team_04_WB.instance_to_wrap.CPU_DAT_O\[9\] _07353_ _07239_ vssd1 vssd1 vccd1
+ vccd1 _07387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11851_ net652 net260 vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _04920_ _06287_ _06288_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__and4bb_2
XANTENNA__12979__B1 net314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ net1285 vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11782_ net758 _05800_ net687 _07267_ _07266_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12443__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13521_ _07743_ _07845_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10733_ _04557_ net635 net550 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__mux2_1
XANTENNA__08742__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ team_04_WB.MEM_SIZE_REG_REG\[30\] net1083 vssd1 vssd1 vccd1 vccd1 _02843_
+ sky130_fd_sc_hd__and2b_1
X_16240_ clknet_leaf_190_wb_clk_i _01909_ _00469_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[213\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input94_A wbs_dat_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ net1552 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[17\] vssd1
+ vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12403_ net519 net600 _07290_ net432 net1897 vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a32o_1
X_13383_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[7\] team_04_WB.MEM_SIZE_REG_REG\[9\]
+ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09072__A1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16171_ clknet_leaf_23_wb_clk_i _01840_ _00400_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[144\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _06135_ net1551 net1022 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09576__S net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15122_ net1246 vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__inv_2
X_12334_ net2204 net499 _07611_ net443 vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
XANTENNA__15875__Q team_04_WB.instance_to_wrap.CPU_DAT_O\[29\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13156__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15053_ net1152 vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12265_ net2396 net505 _07575_ net456 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12903__B1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ net2659 net1070 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__and2_1
X_11216_ net640 _04030_ net360 vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__a21o_1
X_12196_ net2092 net510 _07539_ net458 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12015__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11147_ _06238_ _06245_ net559 vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__mux2_1
XANTENNA__14511__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13459__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14120__A2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15955_ clknet_leaf_72_wb_clk_i _01631_ _00184_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11078_ net572 _06555_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10029_ net591 _04387_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__o21a_1
X_14906_ net1151 vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__inv_2
XANTENNA__12031__A net243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15886_ clknet_leaf_123_wb_clk_i _01563_ _00113_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__dfrtp_1
X_14837_ net1200 vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__inv_2
XANTENNA__13561__S net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__A _05466_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_711 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14768_ net1175 vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16507_ clknet_leaf_101_wb_clk_i _02176_ _00736_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\]
+ sky130_fd_sc_hd__dfrtp_1
X_13719_ _03107_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14699_ net1161 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__inv_2
X_16438_ clknet_leaf_11_wb_clk_i _02107_ _00667_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[411\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13797__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12198__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16369_ clknet_leaf_179_wb_clk_i _02038_ _00598_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13147__B1 net296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11748__C _07216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout305 _07681_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__buf_4
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout316 net317 vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_4
XANTENNA__13736__S net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[609\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__mux2_1
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_4
Xfanout338 net339 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_4
X_17304__1360 vssd1 vssd1 vccd1 vccd1 _17304__1360/HI net1360 sky130_fd_sc_hd__conb_1
Xfanout349 net350 vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__buf_2
XFILLER_0_158_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10920__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__S0 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14111__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _03662_ _05350_ _05351_ _05352_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout281_A _05523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout379_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[34\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[2\]
+ net891 vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10684__A1 team_04_WB.instance_to_wrap.final_design.uart.working_data\[8\]
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ _04232_ _04233_ _04234_ _04235_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04236_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__10684__B2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1190_A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__A _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1288_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08556_ net751 net744 _03726_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__a21oi_4
XANTENNA__13622__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_122_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08487_ _04094_ _04095_ _04096_ _04097_ net784 net800 vssd1 vssd1 vccd1 vccd1 _04098_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12976__A3 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A _03675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout334_X net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1076_X net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10683__X _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12815__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__A1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09396__S net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[749\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[717\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__mux2_1
XANTENNA__08801__A1 _04411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ net617 _05965_ _05620_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or3b_1
XFILLER_0_116_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13138__B1 net295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[236\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[204\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__A team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12050_ net2568 net517 _07478_ net456 vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a22o_1
Xhold370 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] vssd1 vssd1
+ vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[254\] vssd1 vssd1
+ vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _06324_ _06489_ _06322_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__a21oi_1
Xhold392 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\] vssd1 vssd1
+ vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout850 net853 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__clkbuf_4
Xfanout861 net871 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14102__A2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 net873 vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout883 net895 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__clkbuf_4
Xfanout894 net895 vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__buf_2
XANTENNA__12113__B2 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15740_ net1284 vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__inv_2
XANTENNA__10124__B1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_161_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12952_ net230 net2391 net320 vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__mux2_1
Xhold1070 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[643\] vssd1 vssd1
+ vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[876\] vssd1 vssd1
+ vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ net705 _05923_ _07371_ _07372_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__o211a_1
Xhold1092 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[152\] vssd1 vssd1
+ vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ net1282 vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__inv_2
XANTENNA__10675__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _07583_ net342 net390 net2207 vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11690__A net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14622_ net1217 vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__inv_2
X_11834_ net693 _06857_ _07312_ net615 vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12416__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17341_ net1397 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14553_ net1186 vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__inv_2
XFILLER_0_135_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11765_ team_04_WB.instance_to_wrap.CPU_DAT_O\[30\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07253_ sky130_fd_sc_hd__a21o_1
XANTENNA__08715__S1 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_wb_clk_i clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_165_360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13504_ team_04_WB.ADDR_START_VAL_REG\[26\] _02894_ vssd1 vssd1 vccd1 vccd1 _02895_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_155_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10716_ _05473_ net465 vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__nor2_1
X_17272_ team_04_WB.instance_to_wrap.final_design.h_out vssd1 vssd1 vccd1 vccd1 net174
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input97_X net97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11696_ team_04_WB.MEM_SIZE_REG_REG\[26\] _06515_ vssd1 vssd1 vccd1 vccd1 _07185_
+ sky130_fd_sc_hd__xnor2_1
X_14484_ net1163 vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_11_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16223_ clknet_leaf_156_wb_clk_i _01892_ _00452_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[196\]
+ sky130_fd_sc_hd__dfrtp_1
X_13435_ net1082 team_04_WB.MEM_SIZE_REG_REG\[27\] vssd1 vssd1 vccd1 vccd1 _07861_
+ sky130_fd_sc_hd__and2_1
X_10647_ net1054 _06174_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09045__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14506__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13410__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13366_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] team_04_WB.MEM_SIZE_REG_REG\[3\]
+ _07790_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ clknet_leaf_40_wb_clk_i _01823_ _00383_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10578_ team_04_WB.instance_to_wrap.CPU_DAT_O\[7\] net1096 net1054 vssd1 vssd1 vccd1
+ vccd1 _06124_ sky130_fd_sc_hd__and3_1
XANTENNA__11849__B _06729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08063__X _03674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09580__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__B1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15105_ net1188 vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__inv_2
X_12317_ _07320_ net668 vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__and2_1
X_13297_ _06159_ _07719_ _07724_ _07718_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__a32o_1
X_16085_ clknet_leaf_32_wb_clk_i _01754_ _00314_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ net236 net672 vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__and2_1
X_15036_ net1128 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08556__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11865__A net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__B2 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ net248 net647 vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__and2_1
XANTENNA__08308__A0 _03894_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ clknet_leaf_97_wb_clk_i _02656_ _01216_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[960\]
+ sky130_fd_sc_hd__dfrtp_1
X_15938_ clknet_leaf_52_wb_clk_i _01615_ _00165_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10666__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_15869_ clknet_leaf_95_wb_clk_i _01546_ _00096_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10768__X _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _04017_ _04018_ _04019_ _04020_ net823 net741 vssd1 vssd1 vccd1 vccd1 _04021_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_171_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09390_ _04997_ _04998_ _04999_ _05000_ net791 net812 vssd1 vssd1 vccd1 vccd1 _05001_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08385__S net910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12407__A2 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08341_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[250\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[218\]
+ net862 vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11091__A1 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08272_ _03879_ _03880_ _03881_ _03882_ net788 net809 vssd1 vssd1 vccd1 vccd1 _03883_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_15_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_17_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09866__B1_N _05404_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13974__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout496_A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12894__A2 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ACK_I vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07987_ _03512_ net1009 _03596_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout663_A _03633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13990__A _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _03615_ _03622_ _03635_ _03656_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o31a_1
XANTENNA__09198__S1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12646__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10657__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[24\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_09657_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[802\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[770\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_X net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ net751 _03656_ _03726_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__a21oi_2
X_09588_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[419\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[387\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08539_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[182\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[150\]
+ net920 vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10557__C net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ net754 _07027_ _07037_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ _06037_ _06072_ net2658 net1006 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12545__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11481_ net634 _04697_ net358 _06885_ _06968_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__o32a_1
XFILLER_0_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11909__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13220_ net82 team_04_WB.MEM_SIZE_REG_REG\[21\] net982 vssd1 vssd1 vccd1 vccd1 _01683_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10432_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] _06001_
+ _06004_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and3_1
XANTENNA__09122__S1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_150_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12582__A1 _07549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _07585_ net379 net297 net2421 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[8\] _05528_ vssd1
+ vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08043__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ net253 net676 vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_59_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ net233 net2566 net304 vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input57_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _05577_ _05636_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__nand2_1
X_16910_ clknet_leaf_27_wb_clk_i _02579_ _01139_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[883\]
+ sky130_fd_sc_hd__dfrtp_1
X_12033_ _07380_ net685 vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__and2_1
XANTENNA__12334__B2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12885__A2 net345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16841_ clknet_leaf_99_wb_clk_i _02510_ _01070_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[814\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__buf_4
Xfanout691 net692 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__buf_4
X_16772_ clknet_leaf_169_wb_clk_i _02441_ _01001_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13984_ _04583_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__nor2_1
X_15723_ net1294 vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ _07249_ _07663_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nor2_2
XANTENNA__13405__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15654_ net1177 vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12866_ _07566_ net331 net388 net2161 vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ net1284 vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11817_ team_04_WB.instance_to_wrap.CPU_DAT_O\[23\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07298_ sky130_fd_sc_hd__a21o_1
X_15585_ net1131 vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_174_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ net226 net2265 net322 vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_174_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17324_ net1380 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_139_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ net1263 vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__inv_2
X_11748_ _05466_ _06200_ _07216_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17255_ net1315 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
XFILLER_0_154_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14467_ net1250 vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
XANTENNA__09018__B2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _06517_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16206_ clknet_leaf_29_wb_clk_i _01875_ _00435_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\]
+ sky130_fd_sc_hd__dfrtp_1
X_13418_ _07745_ _07837_ _07842_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17186_ clknet_leaf_90_wb_clk_i _02798_ _01415_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_14398_ net1283 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ clknet_leaf_121_wb_clk_i _01806_ _00366_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_13349_ _07773_ _07774_ _07770_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ clknet_leaf_20_wb_clk_i _01737_ _00297_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_07910_ team_04_WB.instance_to_wrap.BUSY_O team_04_WB.EN_VAL_REG vssd1 vssd1 vccd1
+ vccd1 _03524_ sky130_fd_sc_hd__nand2b_1
X_15019_ net1160 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__inv_2
X_08890_ net765 _04500_ _04489_ _04483_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12876__A2 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12203__B net647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12628__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13825__B2 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[100\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[68\]
+ net876 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__mux2_1
XANTENNA__11836__B1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13315__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[550\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[518\]
+ net956 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ _04980_ _04981_ _04982_ _04983_ net793 net813 vssd1 vssd1 vccd1 vccd1 _04984_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13053__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout244_A _07340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08324_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1018\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[986\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08843__S net903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ _03696_ _03754_ _03810_ _03865_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__and4_2
XFILLER_0_7_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12365__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A _07661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08186_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[700\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1039_X net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__S net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15973__Q team_04_WB.ADDR_START_VAL_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__07991__A1 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12316__B2 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__A2 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15809__28 clknet_leaf_56_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13209__B _06140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08091__S1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15705__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__A1 net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12619__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__B2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[224\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[192\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__mux2_1
X_10981_ _06445_ _06453_ _06469_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12720_ net1994 net406 net345 _07427_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _07622_ net489 net410 net1988 vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13044__A2 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ _06415_ _06417_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__xnor2_1
X_15370_ net1112 vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__inv_2
X_12582_ _07549_ net487 net418 net1757 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14321_ net1088 _03479_ _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a21oi_1
X_11533_ net286 _07017_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__or3_1
XANTENNA__10584__A team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08471__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17040_ clknet_leaf_192_wb_clk_i _02709_ _01269_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
X_14252_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[9\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\]
+ _03432_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[11\] vssd1 vssd1
+ vccd1 vccd1 _03436_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__B1 _07455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11399__B net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11464_ _06951_ _06952_ _06950_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__or3b_1
XFILLER_0_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13203_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__nor2_4
XFILLER_0_150_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ net1059 _05996_ net1076 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__mux2_1
X_14183_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] _03393_
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[7\] vssd1 vssd1
+ vccd1 vccd1 _03396_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11395_ net587 _06251_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ _05592_ _05625_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nand2_1
X_13134_ _07568_ net368 net294 net2293 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__a22o_1
X_13065_ net240 net2425 net302 vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__mux2_1
XANTENNA__10318__B1 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ _05759_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__or2_1
XANTENNA__12858__A2 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ net2517 net515 _07461_ net437 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12023__B net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16824_ clknet_leaf_147_wb_clk_i _02493_ _01053_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[797\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08928__S net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09613__A _05223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16755_ clknet_leaf_184_wb_clk_i _02424_ _00984_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09487__A1 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13967_ _04138_ net262 net598 _03317_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11294__A1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ net1262 vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__inv_2
X_12918_ _07620_ net345 net387 net1700 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12491__B1 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16686_ clknet_leaf_26_wb_clk_i _02355_ _00915_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[659\]
+ sky130_fd_sc_hd__dfrtp_1
X_13898_ _03190_ _03274_ _03182_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_17_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15637_ net1178 vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__inv_2
XANTENNA__13035__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ _07547_ net342 net394 net1954 vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09759__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_116 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09334__S1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15568_ net1164 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17307_ net1363 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
X_14519_ net1190 vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__inv_2
XANTENNA__13991__B1 _03330_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15499_ net1161 vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__inv_2
XANTENNA__08041__A_N team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_08040_ net1079 net1028 net1024 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\]
+ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a31o_1
X_17238_ net1404 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_71_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12546__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11349__A2 _06824_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[200\] vssd1 vssd1
+ vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ clknet_leaf_92_wb_clk_i _02781_ _01398_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold914 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[929\] vssd1 vssd1
+ vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[988\] vssd1 vssd1
+ vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[768\] vssd1 vssd1
+ vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09494__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[853\] vssd1 vssd1
+ vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[852\] vssd1 vssd1
+ vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net580 _05167_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold969 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\] vssd1 vssd1
+ vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[687\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[655\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__mux2_1
XANTENNA__12849__A2 net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[240\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[208\]
+ net938 vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11809__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09573__S1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09425_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[422\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[390\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13026__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1270_A net1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout626_A _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08573__S net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[808\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[776\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__mux2_1
XANTENNA__15968__Q team_04_WB.ADDR_START_VAL_REG\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_139_wb_clk_i clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08307_ _03900_ _03906_ _03917_ net717 vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__a22o_2
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09287_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[297\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[265\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[893\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[861\]
+ net877 vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12108__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08169_ net767 _03773_ _03779_ _03761_ _03767_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_127_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10200_ net619 _05803_ _05806_ net280 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_56_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ _06279_ net288 vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _05727_ _05741_ _05726_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_128_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12124__A _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10062_ _03496_ net660 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_145_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ net1229 vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__inv_2
X_13821_ _06840_ net273 vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__nor2_1
XANTENNA__11682__B _07016_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16540_ clknet_leaf_126_wb_clk_i _02209_ _00769_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[513\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11276__A1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13752_ _03122_ _03142_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__or2_1
XANTENNA__12473__B1 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ _06379_ _06448_ _06450_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__a211oi_2
X_12703_ net2146 net404 net326 _07321_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16471_ clknet_leaf_167_wb_clk_i _02140_ _00700_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[444\]
+ sky130_fd_sc_hd__dfrtp_1
X_13683_ team_04_WB.ADDR_START_VAL_REG\[1\] _03073_ vssd1 vssd1 vccd1 vccd1 _03074_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__13017__A2 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ _05084_ _06284_ net659 vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__a21o_1
XANTENNA__13242__X _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09579__S net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ net1236 vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__inv_2
XANTENNA__15170__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ _07605_ net484 net409 net1754 vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11579__A2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15353_ net1245 vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__inv_2
X_12565_ _07532_ net479 net416 net1866 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ net2639 _03467_ net818 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11516_ net567 _06922_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15284_ net1227 vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__inv_2
X_12496_ _07493_ net485 net424 net1646 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__a22o_1
XANTENNA__12528__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ clknet_leaf_159_wb_clk_i _02692_ _01252_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[996\]
+ sky130_fd_sc_hd__dfrtp_1
X_14235_ net2411 _03423_ _03425_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11447_ _06436_ _06903_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_169_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11200__A1 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[1\]
+ _03368_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__and3_1
X_11378_ _06364_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10329_ _05918_ _05921_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[13\]
+ net1075 vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__o2bb2a_1
X_13117_ _07549_ net376 net300 net2043 vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a22o_1
X_14097_ _03518_ _07698_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\] _03516_
+ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__a2bb2o_1
X_13048_ _07509_ net379 net308 net1679 vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__a22o_1
Xfanout1250 net1251 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_4
Xfanout1261 net1297 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__buf_2
XANTENNA__12321__X _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08658__S net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1272 net1273 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_4
Xfanout1283 net1288 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__buf_4
Xfanout1294 net1296 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_1_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16807_ clknet_leaf_166_wb_clk_i _02476_ _01036_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[780\]
+ sky130_fd_sc_hd__dfrtp_1
X_14999_ net1226 vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__inv_2
XFILLER_0_152_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16738_ clknet_leaf_149_wb_clk_i _02407_ _00967_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[711\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__B1 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16669_ clknet_leaf_133_wb_clk_i _02338_ _00898_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[642\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09210_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[234\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[202\]
+ net914 vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__mux2_1
XANTENNA__09489__S net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12216__B1 _07549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09141_ net718 _04751_ _04740_ _04739_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_127_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12209__A _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09072_ net728 _04682_ net713 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_170_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08023_ net760 _03622_ net754 _03631_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__or4_4
XFILLER_0_47_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold700 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[573\] vssd1 vssd1
+ vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10952__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[349\] vssd1 vssd1
+ vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[330\] vssd1 vssd1
+ vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold733 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\] vssd1 vssd1
+ vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[851\] vssd1 vssd1
+ vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold755 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[81\] vssd1 vssd1
+ vccd1 vccd1 net2192 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08294__S1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[308\] vssd1 vssd1
+ vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[472\] vssd1 vssd1
+ vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[891\] vssd1 vssd1
+ vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _04724_ _04727_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__nor2_1
Xhold799 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[967\] vssd1 vssd1
+ vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[431\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[399\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__mux2_1
XANTENNA__13982__B _03308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08856_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[753\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[721\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ net722 _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_140_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout910_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12818__S net324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[807\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[775\]
+ net877 vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__mux2_1
X_10680_ net1763 net1017 net1013 team_04_WB.instance_to_wrap.CPU_DAT_O\[1\] vssd1
+ vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
XANTENNA__09700__B net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12758__A1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\]
+ net890 vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_78_wb_clk_i_A clknet_4_15__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_118_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ net2070 net501 _07619_ net451 vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11981__A2 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ _06246_ _06789_ _06271_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12281_ net2485 net505 _07583_ net453 vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__a22o_1
XANTENNA__12553__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14334__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14020_ _07688_ net1040 _03346_ net1071 net2578 vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_75_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11232_ _06631_ _06634_ net573 vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__mux2_1
XANTENNA__11677__B _07165_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13956__A_N _03807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10581__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ team_04_WB.MEM_SIZE_REG_REG\[26\] _06515_ team_04_WB.MEM_SIZE_REG_REG\[27\]
+ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_112_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_wb_clk_i clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14132__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _05723_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_164_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15971_ clknet_leaf_53_wb_clk_i _01647_ _00200_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_11094_ net634 net546 vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_164_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09234__S0 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _05548_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nand2_1
X_14922_ net1117 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__inv_2
XANTENNA__11497__A1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12694__B1 net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[14\] vssd1 vssd1
+ vccd1 vccd1 net1497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[3\] vssd1
+ vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[3\]
+ vssd1 vssd1 vccd1 vccd1 net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08362__B2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14853_ net1111 vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold93 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[0\]
+ vssd1 vssd1 vccd1 vccd1 net1530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12301__B net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13804_ _03181_ _03190_ _03179_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__a21oi_1
X_14784_ net1213 vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__inv_2
XANTENNA__08114__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ net2350 net517 _07451_ net440 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a22o_1
X_16523_ clknet_leaf_16_wb_clk_i _02192_ _00752_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[496\]
+ sky130_fd_sc_hd__dfrtp_1
X_13735_ net1001 _03125_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10947_ net631 _06433_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14509__A net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16454_ clknet_leaf_17_wb_clk_i _02123_ _00683_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[427\]
+ sky130_fd_sc_hd__dfrtp_1
X_13666_ _03056_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10878_ net635 _06365_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__xor2_2
XFILLER_0_155_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09102__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15405_ net1143 vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__inv_2
XANTENNA__13946__B1 net103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12617_ _07586_ net489 net414 net2308 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a22o_1
X_16385_ clknet_leaf_133_wb_clk_i _02054_ _00614_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[358\]
+ sky130_fd_sc_hd__dfrtp_1
X_13597_ net999 _02987_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__nand2_1
XANTENNA__12029__A _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15336_ net1125 vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__inv_2
XANTENNA__11421__A1 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ net2365 net223 net422 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__mux2_1
XANTENNA__13961__A3 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11972__A2 _07089_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15267_ net1168 vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__inv_2
XANTENNA_2 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net2343 net430 _07652_ net523 vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
XANTENNA__10772__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17006_ clknet_leaf_28_wb_clk_i _02675_ _01235_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[979\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13174__A1 _07610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ _03364_ _03416_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[8\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11587__B _07075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15198_ net1214 vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_state\[1\]
+ sky130_fd_sc_hd__nor2_1
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_120_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09772__S net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14123__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09225__S0 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ net772 _04320_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__or2_1
XANTENNA__15075__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[578\]
+ net892 vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__mux2_1
Xfanout1080 _03523_ vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__clkbuf_2
Xfanout1091 team_04_WB.instance_to_wrap.final_design.VGA_data_control.h_count\[1\]
+ vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__clkbuf_4
X_08641_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[373\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__mux2_1
XANTENNA__12211__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1014\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[982\]
+ net851 vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10947__A net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_112_wb_clk_i_A clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_159_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14138__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout324_A net325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09124_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[301\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08851__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11778__A net653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ _04662_ _04663_ _04664_ _04665_ net786 net806 vssd1 vssd1 vccd1 vccd1 _04666_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__12373__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08006_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1010 _03593_ _03595_ _03590_
+ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_163_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold530 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[864\] vssd1 vssd1
+ vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[353\] vssd1 vssd1
+ vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold552 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\] vssd1 vssd1
+ vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12912__A1 _07614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[75\] vssd1 vssd1
+ vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\] vssd1 vssd1
+ vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold585 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[161\] vssd1 vssd1
+ vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold596 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[610\] vssd1 vssd1
+ vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14114__B1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09957_ _04329_ _04331_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15981__Q team_04_WB.ADDR_START_VAL_REG\[27\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12676__A0 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _04515_ _04516_ _04517_ _04518_ net828 net735 vssd1 vssd1 vccd1 vccd1 _04519_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__11479__A1 _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__S net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _05496_ _05498_ _04359_ _04414_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__o211ai_1
XANTENNA_clkbuf_leaf_151_wb_clk_i_A clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold1230 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[4\] vssd1
+ vssd1 vccd1 vccd1 net2667 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[401\] _03656_ _04449_
+ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__A team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15713__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11850_ _07323_ _07325_ _07326_ net613 vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__o211a_2
XANTENNA__09519__S1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_154_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_154_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12979__A1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10801_ _04584_ _04642_ _06289_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_68_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] net269 net267 vssd1 vssd1 vccd1
+ vccd1 _07267_ sky130_fd_sc_hd__a21o_1
XANTENNA__12548__S net422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13520_ _06681_ net273 vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ net634 _04724_ net546 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08327__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13928__B1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ net1082 team_04_WB.MEM_SIZE_REG_REG\[30\] vssd1 vssd1 vccd1 vccd1 _02842_
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_24_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ net1527 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[18\] vssd1
+ vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a22o_1
X_12402_ net521 net603 _07284_ net433 net1597 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16170_ clknet_leaf_109_wb_clk_i _01839_ _00399_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[143\]
+ sky130_fd_sc_hd__dfrtp_1
X_13382_ _07806_ _07807_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and2_1
XANTENNA_input87_A wbs_dat_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10594_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[2\]
+ _06134_ net1049 vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__mux2_1
XANTENNA__08761__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12600__B1 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ net1272 vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12333_ _07374_ net668 vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__and2_2
XFILLER_0_133_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15052_ net1119 vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12264_ net255 net675 vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_190_wb_clk_i_A clknet_4_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12903__A1 _07605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14003_ net1678 net1069 _03337_ net264 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a22o_1
X_11215_ _04031_ net363 vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__or2_1
X_12195_ net256 net650 vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__and2_1
XANTENNA__14105__B1 _07706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_X net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__X _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ net573 _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__nor2_1
XANTENNA__13459__A2 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12667__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ clknet_leaf_72_wb_clk_i _01630_ _00183_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10531__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11077_ net559 _06560_ _06562_ _06565_ net572 vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08335__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _05572_ _05637_ _05574_ _05571_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__a211o_1
X_14905_ net1241 vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__inv_2
X_15885_ clknet_leaf_124_wb_clk_i _01562_ _00112_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__dfrtp_1
XANTENNA__12031__B net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14836_ net1208 vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__inv_2
XANTENNA__12419__B1 net435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13092__B1 net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14767_ net1143 vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11979_ net692 _07115_ _07437_ net614 vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__o211a_4
XFILLER_0_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16506_ clknet_leaf_38_wb_clk_i _02175_ _00735_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08194__S0 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13718_ _03099_ _03103_ _03106_ team_04_WB.ADDR_START_VAL_REG\[11\] vssd1 vssd1 vccd1
+ vccd1 _03109_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14698_ net1106 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16437_ clknet_leaf_36_wb_clk_i _02106_ _00666_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[410\]
+ sky130_fd_sc_hd__dfrtp_1
X_13649_ net1101 _05526_ net995 _03039_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12198__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16368_ clknet_leaf_192_wb_clk_i _02037_ _00597_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[341\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09694__S0 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15319_ net1229 vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16299_ clknet_leaf_25_wb_clk_i _01968_ _00528_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[272\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_32 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__buf_4
X_09811_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[673\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\]
+ net894 vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__mux2_1
Xfanout317 _07677_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_4
Xfanout328 net332 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__buf_2
Xfanout339 _07667_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_2
XANTENNA__13318__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[416\] _03650_ _03652_
+ _03659_ _03661_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__o311a_1
XANTENNA__09749__S1 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[98\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[66\]
+ net887 vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__mux2_1
XANTENNA__11330__B1 team_04_WB.MEM_SIZE_REG_REG\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_A net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08624_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[948\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[916\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11881__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[15\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11780__B _06185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__A0 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09531__A _05110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ net766 _04165_ _04154_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout441_A net442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12368__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__A3 _07403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12830__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08486_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[55\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[23\]
+ net913 vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__mux2_1
XANTENNA__10396__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13988__A _04752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout706_A net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X net327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[557\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[525\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09038_ _04645_ _04646_ _04647_ _04648_ net789 net811 vssd1 vssd1 vccd1 vccd1 _04649_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12116__B net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold360 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[362\] vssd1 vssd1
+ vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08972__A1_N net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__B1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[316\] vssd1 vssd1
+ vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[355\] vssd1 vssd1
+ vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[438\] vssd1 vssd1
+ vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _06332_ _06482_ _06486_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net843 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
Xfanout851 net853 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12649__B1 net410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout862 net871 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__clkbuf_2
Xfanout873 net874 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__buf_2
Xfanout884 net885 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__buf_4
XANTENNA__12113__A2 net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 net904 vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__buf_2
X_12951_ net232 net2458 net320 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__mux2_1
Xhold1060 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[404\] vssd1 vssd1
+ vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[877\] vssd1 vssd1
+ vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net757 _05925_ _06185_ _04671_ net690 vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__o221a_1
X_15670_ net1282 vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__inv_2
XANTENNA__11872__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[16\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold1082 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[577\] vssd1 vssd1
+ vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08756__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12882_ _07582_ net343 net390 net2102 vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__a22o_1
Xhold1093 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[532\] vssd1 vssd1
+ vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ net1149 vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__inv_2
X_11833_ net704 _05851_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__o21a_1
XANTENNA__13074__A0 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__A team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17340_ net1396 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14552_ net1178 vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__inv_2
XANTENNA__12821__A0 net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11764_ net2094 net527 _07247_ net448 vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_161_Right_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13503_ net996 _02890_ _02893_ _02887_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17271_ net1331 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _05470_ _06201_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_155_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ net1239 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__inv_2
XFILLER_0_165_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11695_ _07170_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16222_ clknet_leaf_143_wb_clk_i _01891_ _00451_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[195\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09587__S net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ net1082 team_04_WB.MEM_SIZE_REG_REG\[27\] vssd1 vssd1 vccd1 vccd1 _07860_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07896__A team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10646_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08491__S net911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output193_A net193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__B1 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ clknet_leaf_177_wb_clk_i _01822_ _00382_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\]
+ sky130_fd_sc_hd__dfrtp_1
X_13365_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] team_04_WB.MEM_SIZE_REG_REG\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nand2_1
XANTENNA__10526__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_51_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10577_ _06123_ net1535 net1021 vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XANTENNA__12307__A _07289_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ net1213 vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ net2197 net499 _07602_ net436 vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a22o_1
X_16084_ clknet_leaf_7_wb_clk_i _01753_ _00313_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_13296_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[1\] team_04_WB.instance_to_wrap.final_design.uart.bits_received\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15035_ net1145 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__inv_2
X_12247_ net2294 net503 _07566_ net443 vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a22o_1
XANTENNA__14522__A net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12888__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__X _04786_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12352__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ net2001 net507 _07530_ net438 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
X_11129_ _06219_ _06221_ net539 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_39_wb_clk_i _02655_ _01215_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[959\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08308__A1 _03918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15937_ clknet_leaf_52_wb_clk_i _01614_ _00164_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11312__A0 _03891_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__A1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__A2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15868_ clknet_leaf_98_wb_clk_i _01545_ _00095_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_14819_ net1170 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11092__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12812__A0 _07385_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[58\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[26\]
+ net867 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08271_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[955\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[923\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__B team_04_WB.MEM_SIZE_REG_REG\[18\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12040__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__A net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12591__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12879__B1 net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_1066 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout391_A _07673_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_A net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ _03512_ net1009 _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_35_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13990__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ net768 _05335_ _05324_ _05323_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__o2bb2a_4
XTAP_TAPCELL_ROW_87_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11854__A1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__A2 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[866\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[834\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08576__S net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_91 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ net766 _04217_ _04206_ _04205_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__o2bb2a_4
XANTENNA_fanout823_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[483\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[451\]
+ net957 vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout444_X net444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1186_X net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10409__A2 net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__A0 _07327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08538_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[246\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[214\]
+ net919 vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _04074_ _04079_ net721 vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[0\]
+ _06051_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_133_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11480_ _04668_ _04697_ net361 vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__a21o_1
XANTENNA__14020__A2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[4\] _06009_
+ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ _07584_ net376 net296 net1970 vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a22o_1
XANTENNA__12582__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] _05950_ net1076
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12101_ net2228 net352 _07505_ net442 vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
XANTENNA__08043__C net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10293_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[17\] _05889_ net1075
+ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ net261 net2449 net304 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__mux2_1
XANTENNA__12334__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ net2417 net516 _07469_ net449 vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
Xhold190 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[165\] vssd1 vssd1
+ vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ clknet_leaf_116_wb_clk_i _02509_ _01069_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout670 _07589_ vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_4
XANTENNA__11972__Y _07432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout681 net685 vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__clkbuf_8
Xfanout692 _06187_ vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__clkbuf_4
X_16771_ clknet_leaf_125_wb_clk_i _02440_ _01000_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[744\]
+ sky130_fd_sc_hd__dfrtp_1
X_13983_ _07344_ _03308_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__or2_1
X_15722_ net1296 vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ net246 net2589 net318 vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15653_ net1177 vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__inv_2
XANTENNA__13405__B team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ _07565_ net328 net388 net1893 vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__a22o_1
XANTENNA__13047__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output206_A net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08149__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13598__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14604_ net1287 vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ net758 _05837_ net697 _04113_ net693 vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__a221o_1
X_15584_ net1153 vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ net227 net2370 net323 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_174_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ net1379 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_133_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_174_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_174_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11747_ _06200_ net271 vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17254_ net1314 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_126_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14466_ net1272 vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__inv_2
X_11678_ team_04_WB.MEM_SIZE_REG_REG\[28\] _06516_ vssd1 vssd1 vccd1 vccd1 _07167_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10764__B _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ clknet_leaf_42_wb_clk_i _01874_ _00434_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[178\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13417_ _07745_ _07842_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10629_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[13\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[12\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[15\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[14\]
+ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__or4_1
X_17185_ clknet_leaf_90_wb_clk_i _02797_ _01414_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14397_ net1287 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12037__A net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xmax_cap804 _03551_ vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
XFILLER_0_113_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12573__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ clknet_leaf_113_wb_clk_i _01805_ _00365_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[6\] team_04_WB.MEM_SIZE_REG_REG\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11876__A net656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15348__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ clknet_leaf_118_wb_clk_i _01736_ _00296_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_13279_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\] _07710_ _05525_
+ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__mux2_1
XANTENNA__09726__B1 _03656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ net1116 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16969_ clknet_leaf_100_wb_clk_i _02638_ _01198_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[942\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08388__S0 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[164\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[132\]
+ net879 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__mux2_1
XANTENNA__13155__X _07684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08396__S net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__X _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_215 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09441_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[614\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[582\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13038__B1 net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09372_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[423\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[391\]
+ net945 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_83 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08323_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[794\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12261__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10811__A2 _06291_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ _03834_ _03861_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09020__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13210__A0 net93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08185_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[764\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[732\]
+ net879 vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout404_A _07664_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12564__A2 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13761__B2 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__B1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12381__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12316__A2 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09256__A net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11524__A0 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13209__C _06145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09690__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11792__Y _07277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07969_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1023\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[991\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout940_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout659_X net659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[32\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[0\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__mux2_1
XANTENNA__11827__A1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _06357_ _06463_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__or3_1
XANTENNA__12410__A net651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09639_ net664 _05248_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a21o_1
XANTENNA__13029__B1 net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12650_ _07621_ net489 net410 net1948 vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11601_ net708 _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12581_ _07548_ net490 net418 net1796 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__a22o_1
XANTENNA__14337__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14320_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[31\]
+ _03357_ _03471_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[30\]
+ net1087 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_262 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11532_ _06278_ _07015_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10584__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ net2620 _03433_ _03435_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__B2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11463_ _04867_ _06248_ net362 _04866_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__a22o_1
X_13202_ team_04_WB.instance_to_wrap.wb_manage.curr_state\[0\] _07695_ _07698_ vssd1
+ vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__and3_1
X_10414_ net1059 net283 _05993_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22oi_1
XANTENNA__12555__A2 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ net2666 _03393_ _03395_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[6\]
+ sky130_fd_sc_hd__a21oi_1
X_11394_ _06378_ _06882_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13133_ _07567_ net367 net294 net2077 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__a22o_1
XANTENNA__15168__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ net2655 net1057 _05932_ _05935_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13064_ net242 net2529 net302 vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__mux2_1
XANTENNA__10318__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ _05692_ _05758_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_167_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ net246 net680 vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__and2_1
XANTENNA__14800__A net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13268__A0 net99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16823_ clknet_leaf_175_wb_clk_i _02492_ _01052_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11530__A3 _06272_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11818__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16754_ clknet_leaf_6_wb_clk_i _02423_ _00983_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[727\]
+ sky130_fd_sc_hd__dfrtp_1
X_13966_ net151 net1065 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15705_ net1258 vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__inv_2
X_12917_ _07619_ net341 net386 net2341 vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__a22o_1
XANTENNA__11294__A2 _06781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12491__A1 _07488_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16685_ clknet_leaf_32_wb_clk_i _02354_ _00914_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[658\]
+ sky130_fd_sc_hd__dfrtp_1
X_13897_ _03148_ _03192_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_17_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15636_ net1178 vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__inv_2
XFILLER_0_159_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12848_ _07546_ net343 net394 net1793 vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__a22o_1
XANTENNA__08944__S net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15567_ net1195 vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12243__B2 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ _07506_ net330 net396 net2109 vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a22o_1
XANTENNA__10775__A _03721_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12319__X _07604_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17306_ net1362 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
X_14518_ net1190 vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__inv_2
XANTENNA__10254__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08542__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15498_ net1107 vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__inv_2
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14449_ net1276 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__inv_2
X_17237_ net1403 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_141_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17168_ clknet_leaf_93_wb_clk_i _02780_ _01397_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold904 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[292\] vssd1 vssd1
+ vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold915 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[479\] vssd1 vssd1
+ vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[664\] vssd1 vssd1
+ vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16119_ clknet_leaf_161_wb_clk_i _01788_ _00348_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold937 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[282\] vssd1 vssd1
+ vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_4_4__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold948 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[906\] vssd1 vssd1
+ vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17099_ clknet_leaf_76_wb_clk_i _02734_ _01328_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_09990_ net580 _05167_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__or2_1
Xhold959 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[845\] vssd1 vssd1
+ vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08941_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[751\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[719\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12989__X _07678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08872_ net772 _04482_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_32_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13259__A0 net77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11809__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12823__C_N net650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__S net900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout354_A net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08781__S0 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[486\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[454\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08854__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09355_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[840\]
+ net900 vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__mux2_1
XANTENNA__11037__A2 net581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12376__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout521_A net522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ _03911_ _03916_ net722 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_A clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12785__A2 net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09286_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[361\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[329\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08237_ net730 _03847_ net714 vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__o21a_1
XANTENNA__13996__A _04918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_wb_clk_i clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_179_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__09685__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ net780 _03778_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08099_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[894\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\]
+ net942 vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10130_ _05730_ _05740_ _05729_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _03496_ net660 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13820_ _03209_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_162_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ _03132_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__nand2_1
X_10963_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__inv_2
XANTENNA__12473__A1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12702_ net2184 net404 net326 _07314_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16470_ clknet_leaf_11_wb_clk_i _02139_ _00699_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[443\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13682_ net1001 _03071_ _03072_ _03069_ _03070_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a32o_1
XANTENNA__08764__S net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10894_ _06381_ _06382_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15421_ net1153 vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12633_ _07604_ net484 net409 net1630 vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15352_ net1204 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12776__A2 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13973__A1 _04243_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12564_ _07531_ net481 net416 net1684 vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14303_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\] _03467_
+ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11515_ net555 _06960_ _06961_ _07003_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15283_ net1231 vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ _07492_ net481 net424 net1955 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17022_ clknet_leaf_116_wb_clk_i _02691_ _01251_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[995\]
+ sky130_fd_sc_hd__dfrtp_1
X_14234_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[4\] _03423_ net820
+ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_117_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input72_X net72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11446_ team_04_WB.MEM_SIZE_REG_REG\[10\] _06504_ vssd1 vssd1 vccd1 vccd1 _06935_
+ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14165_ _03383_ _03384_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.v_next_count\[0\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_169_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__S net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11200__A2 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_890 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11377_ _06367_ _06865_ _06366_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13116_ _07548_ net378 net300 net1952 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a22o_1
X_10328_ net282 _05920_ net1057 vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a21oi_1
X_14096_ net1530 _06138_ net1034 vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__mux2_1
X_13047_ _07508_ net380 net309 net2038 vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__a22o_1
X_10259_ net280 _05857_ net1056 vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21oi_1
Xfanout1240 net1242 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__buf_2
XANTENNA__09624__A net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12700__A2 net404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1251 net1252 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__buf_4
Xfanout1262 net1264 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10172__C1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1273 net1279 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__buf_4
Xfanout1284 net1288 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_1_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_53_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1295 net1296 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__buf_4
X_16806_ clknet_leaf_20_wb_clk_i _02475_ _01035_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[779\]
+ sky130_fd_sc_hd__dfrtp_1
X_14998_ net1228 vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__inv_2
XFILLER_0_163_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16737_ clknet_leaf_135_wb_clk_i _02406_ _00966_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__A1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A2 _06750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _05338_ net710 _03307_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or3_4
XFILLER_0_163_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_102_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08674__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16668_ clknet_leaf_127_wb_clk_i _02337_ _00897_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08527__X _04138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13008__A3 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15619_ net1170 vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12216__B2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16599_ clknet_leaf_174_wb_clk_i _02268_ _00828_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[572\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10227__B1 net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12767__A2 net329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09140_ _04745_ _04750_ net730 vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_wb_clk_i clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12209__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_62_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09071_ _04678_ _04679_ _04680_ _04681_ net829 net736 vssd1 vssd1 vccd1 vccd1 _04682_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12924__S net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08840__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08022_ net757 _03623_ net708 net705 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__and4_1
XANTENNA__12519__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[521\] vssd1 vssd1
+ vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08703__A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold712 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[332\] vssd1 vssd1
+ vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1015\] vssd1 vssd1
+ vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold734 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[879\] vssd1 vssd1
+ vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[947\] vssd1 vssd1
+ vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold756 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[209\] vssd1 vssd1
+ vccd1 vccd1 net2193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[812\] vssd1 vssd1
+ vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[855\] vssd1 vssd1
+ vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05583_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold789 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[873\] vssd1 vssd1
+ vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[463\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1011_A _03547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08849__S net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09699__A2 _05307_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08855_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[561\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[529\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout471_A _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout569_A _05251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08786_ _04393_ _04394_ _04395_ _04396_ net827 net743 vssd1 vssd1 vccd1 vccd1 _04397_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_140_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09821__X _05432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_A net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__B2 net520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A team_04_WB.instance_to_wrap.CPU_DAT_O\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[871\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[839\]
+ net884 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A net904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12758__A2 net334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09338_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[104\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[72\]
+ net893 vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__mux2_1
XANTENNA__13955__A1 _03860_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ net779 _04879_ net761 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ _05475_ _06788_ net563 vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12280_ net224 net674 vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout893_X net893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_180_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13183__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ _06246_ _06632_ _06271_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12391__A0 _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__C net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _06638_ _06650_ net464 _06630_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_112_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10113_ _03724_ _04002_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_164_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15970_ clknet_leaf_50_wb_clk_i _01646_ _00199_ vssd1 vssd1 vccd1 vccd1 team_04_WB.ADDR_START_VAL_REG\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14350__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12143__A0 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _06580_ _06581_ net539 vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09234__S1 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input32_A DAT_I[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ net643 _03836_ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21o_1
X_14921_ net1133 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__inv_2
Xhold50 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[6\] vssd1
+ vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_76_wb_clk_i clknet_4_13__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold61 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[4\] vssd1
+ vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 _02763_ vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[9\] vssd1 vssd1
+ vccd1 vccd1 net1520 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ net1169 vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__inv_2
Xhold94 net166 vssd1 vssd1 vccd1 vccd1 net1531 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _03148_ _03170_ _03193_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__or3_2
X_14783_ net1241 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11995_ net212 net682 vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__and2_1
X_13734_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[9\] net1045 _03124_
+ net1093 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12997__A2 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16522_ clknet_leaf_164_wb_clk_i _02191_ _00751_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[495\]
+ sky130_fd_sc_hd__dfrtp_1
X_10946_ net631 _06433_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_119_Left_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13665_ _03054_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__or2_1
X_16453_ clknet_leaf_20_wb_clk_i _02122_ _00682_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[426\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10529__S net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ net635 _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12749__A2 net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _07585_ net489 net414 net2377 vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a22o_1
X_15404_ net1120 vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__inv_2
XANTENNA__13946__B2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16384_ clknet_leaf_135_wb_clk_i _02053_ _00613_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_716 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13596_ net995 _02984_ _02986_ _07691_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12029__B net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ net1142 vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__inv_2
X_12547_ net2299 net234 net422 vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__mux2_1
XANTENNA__11421__A2 _04724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14525__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ net1219 vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__inv_2
XANTENNA__08082__X _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ net607 net232 net682 vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__and3_1
XANTENNA_3 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ net1973 _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.vga.h_next_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_17005_ clknet_leaf_41_wb_clk_i _02674_ _01234_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[978\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13174__A2 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11429_ net755 _06915_ _06917_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__and3_1
XANTENNA__12045__A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15197_ net1154 vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__A0 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14148_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] _03359_
+ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\] vssd1 vssd1 vccd1
+ vccd1 _03369_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12921__A2 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__A1 net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11884__A net655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ net1481 _06104_ net1033 vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__mux2_1
XANTENNA__12134__A0 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09225__S1 net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__A2 _06427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13882__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1070 net1073 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__buf_2
Xfanout1081 _03515_ vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__buf_4
X_08640_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[437\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[405\]
+ net906 vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1092 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\] vssd1
+ vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_2
XANTENNA__11890__Y _07362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08571_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[822\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[790\]
+ net851 vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__mux2_1
XANTENNA__12437__B2 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12988__A2 _07668_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13323__B team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17155__1298 vssd1 vssd1 vccd1 vccd1 _17155__1298/HI net1298 sky130_fd_sc_hd__conb_1
XFILLER_0_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17283__1339 vssd1 vssd1 vccd1 vccd1 _17283__1339/HI net1339 sky130_fd_sc_hd__conb_1
XANTENNA__09161__S0 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[365\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[333\]
+ net898 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__mux2_1
XANTENNA__12654__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout317_A _07677_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[684\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[652\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__mux2_1
XANTENNA__11778__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] net1009 _03593_ _03595_ _03590_
+ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13165__A2 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold520 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\] vssd1 vssd1
+ vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12373__A0 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold531 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1000\] vssd1 vssd1
+ vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold542 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[888\] vssd1 vssd1
+ vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_173 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12912__A2 net330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\] vssd1 vssd1
+ vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[887\] vssd1 vssd1
+ vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__C1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold575 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[126\] vssd1 vssd1
+ vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[957\] vssd1 vssd1
+ vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14114__A1 team_04_WB.MEM_SIZE_REG_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout686_A net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold597 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[881\] vssd1 vssd1
+ vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14114__B2 team_04_WB.ADDR_START_VAL_REG\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ net639 _04219_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_70_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08907_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[816\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[784\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_1
X_09887_ _04475_ _04476_ _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13873__B1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1220 team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[7\] vssd1 vssd1
+ vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout853_A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_X net474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1231 team_04_WB.instance_to_wrap.final_design.uart.working_data\[7\] vssd1 vssd1
+ vccd1 vccd1 net2668 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10687__B1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _03505_ net1008 net1007 _03658_ _03660_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__a311o_1
XPHY_EDGE_ROW_142_Right_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10697__X _06186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[754\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[722\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ _04697_ _04753_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11780_ _03783_ _06185_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_3__f_wb_clk_i_A clknet_3_1_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10731_ _06218_ _06219_ net539 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _07727_ _07870_ _07875_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_24_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10662_ net1533 net1016 net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[19\] vssd1
+ vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11939__B1 net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12401_ net2191 net433 _07629_ net521 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_123_wb_clk_i clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] team_04_WB.MEM_SIZE_REG_REG\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__or2_1
X_10593_ team_04_WB.instance_to_wrap.CPU_DAT_O\[2\] net1096 net1051 vssd1 vssd1 vccd1
+ vccd1 _06134_ sky130_fd_sc_hd__and3_1
XANTENNA__14345__A net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__A _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15120_ net1163 vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ net2492 net502 _07610_ net456 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13156__A2 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15051_ net1160 vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__inv_2
X_12263_ net2325 net506 _07574_ net459 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14002_ _05029_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nor2_1
X_11214_ net571 _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__nand2_1
X_12194_ net2171 net510 _07538_ net451 vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
X_11145_ _06223_ _06232_ net560 vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input35_X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15953_ net1407 _01629_ _00181_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_11076_ net536 _06564_ net559 vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__o21ai_1
X_10027_ _05572_ _05637_ _05574_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__a21o_1
X_14904_ net1205 vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__inv_2
X_15884_ clknet_leaf_123_wb_clk_i _01561_ _00111_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ net1231 vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__inv_2
XANTENNA__12419__A1 net525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13616__B1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A2 _07150_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_127_Left_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11978_ _07398_ _07436_ _07435_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__a21o_1
X_14766_ net1200 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__inv_2
X_16505_ clknet_leaf_178_wb_clk_i _02174_ _00734_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08194__S1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__inv_2
XFILLER_0_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929_ _06415_ _06416_ _06403_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__a21o_1
X_14697_ net1132 vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16436_ clknet_leaf_8_wb_clk_i _02105_ _00665_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[409\]
+ sky130_fd_sc_hd__dfrtp_1
X_13648_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\] _03026_ vssd1
+ vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__nor2_1
XANTENNA__08952__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13579_ _02958_ _02968_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nand2_1
X_16367_ clknet_leaf_187_wb_clk_i _02036_ _00596_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[340\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10783__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09694__S1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_974 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15318_ net1222 vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__inv_2
X_16298_ clknet_leaf_164_wb_clk_i _01967_ _00527_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08253__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_136_Left_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13147__A2 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_44 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15249_ net1273 vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09783__S net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire275_X net275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[737\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\]
+ net893 vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__mux2_1
Xfanout307 _07680_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_4
XANTENNA__12062__X _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout318 net319 vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__buf_6
Xfanout329 net331 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_4
X_09741_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[384\] _03654_ _03655_
+ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__or3_1
XANTENNA__10669__B1 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _03640_ net703 _05277_ _05281_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_145_Left_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08623_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1012\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[980\]
+ net841 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08709__S0 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _04159_ _04164_ net771 vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09531__B net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14280__B1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[119\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[87\]
+ net912 vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout434_A _07625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09134__S0 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12384__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout222_X net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12594__B1 net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[621\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[589\]
+ net949 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09037_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[428\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[396\]
+ net940 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__mux2_1
XANTENNA__13138__A2 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15789__8 clknet_leaf_68_wb_clk_i vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__inv_2
Xhold350 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[173\] vssd1 vssd1
+ vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[703\] vssd1 vssd1
+ vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 net123 vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[245\] vssd1 vssd1
+ vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[499\] vssd1 vssd1
+ vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout830 net838 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout841 net843 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__buf_4
Xfanout852 net853 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__clkbuf_4
X_09939_ net644 _03783_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nand2_1
XANTENNA__08102__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12649__A1 _07620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net871 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__clkbuf_4
Xfanout874 net904 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_2
Xfanout885 net889 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_4
XANTENNA__09514__A1 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ net223 net2246 net320 vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__mux2_1
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11857__C1 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1050 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[0\] vssd1
+ vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ net687 _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
XANTENNA__09281__X _04892_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[269\] vssd1 vssd1
+ vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\] vssd1 vssd1
+ vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
X_12881_ _07581_ net343 net390 net2056 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a22o_1
Xhold1083 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[705\] vssd1 vssd1
+ vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10868__A net636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[862\] vssd1 vssd1
+ vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_107_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ net686 _07310_ _07309_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ net1126 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__inv_2
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_159_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_159_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10587__B net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14551_ net1178 vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__inv_2
XANTENNA__09373__S0 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11763_ _06198_ net611 vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11624__A2 _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ net996 _02892_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__nand2_1
X_10714_ _05470_ _06201_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nor2_1
X_17270_ net1330 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_155_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ net1159 vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__inv_2
X_11694_ net706 _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_165_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13433_ _07858_ _07729_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__and2b_1
X_16221_ clknet_leaf_131_wb_clk_i _01890_ _00450_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[194\]
+ sky130_fd_sc_hd__dfrtp_1
X_10645_ team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[1\] net1098
+ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__or2_2
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12585__B1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_172_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16152_ clknet_leaf_149_wb_clk_i _01821_ _00381_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[125\]
+ sky130_fd_sc_hd__dfrtp_1
X_13364_ _07786_ _07789_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10576_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[8\]
+ _06122_ net1048 vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12307__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11986__X _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ net237 net668 vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__and2_1
XANTENNA__13129__A2 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15103_ net1270 vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16083_ clknet_leaf_188_wb_clk_i _01752_ _00312_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_13295_ team_04_WB.instance_to_wrap.final_design.uart.bits_received\[2\] _07718_
+ _07719_ _07723_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15034_ net1153 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__inv_2
XANTENNA__08005__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12246_ net248 net672 vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_91_wb_clk_i clknet_4_12__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__08556__A2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_47 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ net239 net647 vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_20_wb_clk_i clknet_4_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12323__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__S net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11128_ _06616_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__inv_2
X_16985_ clknet_leaf_151_wb_clk_i _02654_ _01214_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[958\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17282__1338 vssd1 vssd1 vccd1 vccd1 _17282__1338/HI net1338 sky130_fd_sc_hd__conb_1
X_15936_ clknet_leaf_57_wb_clk_i _01613_ _00163_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__dfrtp_1
X_11059_ net639 net543 vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11312__A1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire235_A _07408_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15867_ clknet_leaf_95_wb_clk_i _01544_ _00094_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.CPU_DAT_O\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10778__A net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818_ net1255 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09269__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__S1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14749_ net1149 vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__inv_2
XFILLER_0_171_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09778__S net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[1019\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[987\]
+ net927 vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08682__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10784__Y _06273_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_2__f_wb_clk_i_X clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16419_ clknet_leaf_118_wb_clk_i _02088_ _00648_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[392\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12057__X _07482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12576__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12040__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__B net649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12932__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11226__S1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09744__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07985_ net1079 net1028 net1024 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__a31oi_2
XANTENNA_fanout384_A _07674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _05329_ _05334_ net776 vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__mux2_1
XANTENNA__08857__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13990__C _03325_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__C1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12500__B1 net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__A net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[930\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[898\]
+ net959 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__mux2_1
XANTENNA__12379__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A net1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _04211_ _04216_ net770 vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout649_A _07520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_171_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[291\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[259\]
+ net948 vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08537_ net771 _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout816_A net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__S net892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10814__B1 _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _04075_ _04076_ _04077_ _04078_ net825 net742 vssd1 vssd1 vccd1 vccd1 _04079_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_61_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ net720 _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout604_X net604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__A net652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12567__B1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__S1 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] _06002_
+ _06005_ _06007_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10361_ _05948_ _05949_ net282 vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__mux2_1
XANTENNA__11790__A1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12100_ net254 net677 vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__and2_2
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ net249 net2474 net305 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__mux2_1
XANTENNA__08043__D net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10292_ net278 _05888_ _05886_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__o21a_1
XANTENNA__10870__B _05463_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12031_ net243 net681 vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__and2_1
XANTENNA__10362__S net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[112\] vssd1 vssd1
+ vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[0\] vssd1 vssd1
+ vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10345__A2 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11982__A team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout671 _07589_ vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__buf_2
X_16770_ clknet_leaf_149_wb_clk_i _02439_ _00999_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[743\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout682 net684 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__buf_4
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__buf_4
XANTENNA__08767__S net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13982_ _07344_ _03308_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15721_ net1294 vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__inv_2
XANTENNA__09594__S0 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ net236 net2532 net318 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_126_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15652_ net1177 vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12864_ _07564_ net329 net388 net2220 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a22o_1
X_14603_ net1287 vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08149__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ net2346 net526 net440 _07296_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12795_ net217 net2554 net322 vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__mux2_1
X_15583_ net1270 vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__inv_2
XFILLER_0_157_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_174_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ net1378 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__09598__S net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ net266 vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__inv_2
X_14534_ net1292 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_174_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17253_ net1313 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_12_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14465_ net1285 vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__inv_2
X_11677_ net707 _07165_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__or2_1
XANTENNA__10537__S net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12558__B1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ clknet_leaf_107_wb_clk_i _01873_ _00433_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[177\]
+ sky130_fd_sc_hd__dfrtp_1
X_13416_ _07741_ _07841_ _07744_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_141_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10628_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[29\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[28\]
+ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[31\] team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[30\]
+ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__or4_1
X_17184_ clknet_leaf_87_wb_clk_i _02796_ _01413_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_14396_ net1255 vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12022__A2 net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12037__B net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13347_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[5\] team_04_WB.MEM_SIZE_REG_REG\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16135_ clknet_leaf_24_wb_clk_i _01804_ _00364_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10559_ _06111_ net1576 net1020 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_4_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11781__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[28\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13278_ net617 _07434_ _07709_ _05615_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16066_ clknet_leaf_144_wb_clk_i _01735_ _00295_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11876__B net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08531__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10780__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12229_ net2388 net504 _07557_ net448 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__a22o_1
X_15017_ net1132 vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__inv_2
XANTENNA__12053__A net228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12730__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15364__A net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08677__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16968_ clknet_leaf_114_wb_clk_i _02637_ _01197_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[941\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12089__A2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15919_ clknet_leaf_73_wb_clk_i _01596_ _00146_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__dfrtp_1
XANTENNA__11297__B1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08388__S1 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11836__A2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ clknet_leaf_124_wb_clk_i _02568_ _01128_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[872\]
+ sky130_fd_sc_hd__dfrtp_1
X_09440_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[678\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[646\]
+ net953 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[487\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[455\]
+ net944 vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_474 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12927__S net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12797__A0 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_95 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08322_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[890\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[858\]
+ net928 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_58_wb_clk_i_A clknet_4_7__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12261__A2 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09301__S net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ net643 _03861_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12228__A net211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08184_ net727 _03794_ net714 vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12662__S net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout599_A _03309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A3 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A1 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12721__B1 net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout766_A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[831\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[799\]
+ net932 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
XANTENNA__08587__S net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[96\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[64\]
+ net969 vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[5\] vssd1
+ vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout933_A net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_wb_clk_i_A clknet_4_14__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12410__B net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09638_ net664 _05223_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_168_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09569_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[869\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[837\]
+ net886 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12788__B1 net398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _06205_ _07083_ _07088_ _07079_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a31o_2
XFILLER_0_155_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _07547_ net490 net418 net1601 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09653__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09211__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ net589 _05030_ net358 _07018_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__o311a_1
XFILLER_0_147_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10584__C net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14250_ team_04_WB.instance_to_wrap.final_design.uart.BAUD_counter\[10\] _03433_
+ net820 vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _06887_ _06946_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12004__A2 net516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17281__1337 vssd1 vssd1 vccd1 vccd1 _17281__1337/HI net1337 sky130_fd_sc_hd__conb_1
X_13201_ _05338_ _07235_ net710 vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ net617 _05994_ net283 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__a21oi_1
X_14181_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[6\] _03393_
+ _03373_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ _06373_ _06864_ _06370_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__a21o_1
XANTENNA__10881__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14353__A net1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _07566_ net371 net294 net1918 vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__a22o_1
XANTENNA__12960__B1 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10344_ net279 _05934_ net1076 vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_78_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input62_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13063_ net226 net2564 net302 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__mux2_1
X_10275_ _05571_ _05638_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11515__A1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08916__C1 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ net2552 net515 _07460_ net436 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XANTENNA__12712__B1 net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_167_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08392__B1 _03725_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16822_ clknet_leaf_12_wb_clk_i _02491_ _01051_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12160__X _07521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout490 net491 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09182__A net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16753_ clknet_leaf_172_wb_clk_i _02422_ _00982_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[726\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11818__A2 _07298_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ _04081_ net262 net598 _03316_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a31o_1
X_15704_ net1257 vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__inv_2
X_12916_ _07618_ net342 net386 net2179 vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10121__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16684_ clknet_leaf_110_wb_clk_i _02353_ _00913_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[657\]
+ sky130_fd_sc_hd__dfrtp_1
X_13896_ _03270_ _03273_ net1992 net1067 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_150_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12491__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09910__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ net1178 vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14312__S0 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12847_ _07545_ net347 net395 net1752 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a22o_1
XANTENNA__14528__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12779__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12243__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15566_ net1197 vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12778_ _07505_ net337 net397 net1898 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
XANTENNA__09121__S net896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10775__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17305_ net1361 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__10254__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__A0 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517_ net1192 vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08542__S1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11729_ _06625_ _06626_ _06656_ _07184_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__a211o_1
XANTENNA__13991__A2 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15497_ net1134 vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17236_ net1402 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
X_14448_ net1276 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17167_ clknet_leaf_93_wb_clk_i _02779_ _01396_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10791__A _05464_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold905 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[660\] vssd1 vssd1
+ vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
X_14379_ net1439 vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11754__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12951__A0 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold916 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[156\] vssd1 vssd1
+ vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold927 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[264\] vssd1 vssd1
+ vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ clknet_leaf_14_wb_clk_i _01787_ _00347_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[984\] vssd1 vssd1
+ vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
X_17098_ clknet_leaf_75_wb_clk_i _02733_ _01327_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold949 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[665\] vssd1 vssd1
+ vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08261__A net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16049_ clknet_leaf_184_wb_clk_i _01718_ _00278_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08940_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[559\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[527\]
+ net947 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__mux2_1
XANTENNA__12703__B1 net326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09175__A2 _03644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_131_wb_clk_i_A clknet_4_10__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08871_ _04478_ _04479_ _04480_ _04481_ net789 net811 vssd1 vssd1 vccd1 vccd1 _04482_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_32_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13607__A _07685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10730__S net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13259__A1 team_04_WB.ADDR_START_VAL_REG\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13326__B team_04_WB.MEM_SIZE_REG_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__S net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__B net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__S0 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[294\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[262\]
+ net954 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10493__A1 team_04_WB.instance_to_wrap.final_design.VGA_adr\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08781__S1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__S net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout347_A net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09354_ _04961_ _04962_ _04963_ _04964_ net836 net737 vssd1 vssd1 vccd1 vccd1 _04965_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_164_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09031__S net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ _03912_ _03913_ _03914_ _03915_ net828 net743 vssd1 vssd1 vccd1 vccd1 _03916_
+ sky130_fd_sc_hd__mux4_1
X_09285_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[393\]
+ net857 vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1256_A net1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08236_ _03843_ _03844_ _03845_ _03846_ net831 net737 vssd1 vssd1 vccd1 vccd1 _03847_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08870__S net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13996__B net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11797__A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08167_ _03774_ _03775_ _03776_ _03777_ net791 net812 vssd1 vssd1 vccd1 vccd1 _03778_
+ sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_170_wb_clk_i_A clknet_4_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1044_X net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12942__A0 _07368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ net779 _03708_ net763 vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_56_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout883_A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10206__A net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14901__A net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_148_wb_clk_i clknet_4_8__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_148_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_10060_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[27\] _03894_ vssd1
+ vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_73_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_145_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_167_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_145_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10640__S _06173_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09206__S net914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_162_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15732__A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ team_04_WB.ADDR_START_VAL_REG\[8\] _03139_ vssd1 vssd1 vccd1 vccd1 _03141_
+ sky130_fd_sc_hd__xor2_1
X_10962_ _06362_ _06366_ _06363_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__o21bai_1
XANTENNA__08221__S0 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12473__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A3 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ net2065 net404 net329 _07308_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13681_ team_04_WB.MEM_SIZE_REG_REG\[1\] net1081 net1046 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__o22a_1
X_10893_ _04947_ _06380_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nand2_1
XANTENNA__14348__A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15420_ net1145 vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__inv_2
X_12632_ _07603_ net479 net408 net1953 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__B2 _05525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15351_ net1229 vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ _07530_ net480 net416 net1721 vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13973__A2 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11984__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__10787__A2 _06269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14302_ _03467_ net818 _03466_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__and3b_1
XFILLER_0_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11514_ net563 _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__and2_1
XFILLER_0_163_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09729__X _05340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08780__S net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ _07491_ net479 net424 net1854 vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
X_15282_ net1244 vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ clknet_leaf_131_wb_clk_i _02690_ _01250_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[994\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13186__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ _06509_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__and2_1
X_14233_ _03423_ _03424_ net819 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08288__S0 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11736__A1 _06816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12933__A0 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_169_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14164_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.v_count\[0\] _03368_
+ _03382_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_169_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11376_ _06373_ _06377_ _06864_ _06449_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12315__B net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ _05532_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__nor2_1
X_13115_ _07547_ net378 net300 net2046 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14095_ net1505 _06136_ net1034 vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__mux2_1
X_13046_ _07507_ net372 net306 net1883 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__a22o_1
X_10258_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_38 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1230 net1253 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__clkbuf_4
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__buf_4
XFILLER_0_79_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ _05551_ _05652_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12331__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1252 net1253 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_2
Xfanout1263 net1264 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_4
Xfanout1274 net1279 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__buf_4
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__buf_4
X_16805_ clknet_leaf_185_wb_clk_i _02474_ _01034_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[778\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1296 net1297 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
XANTENNA__08117__B1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ net1211 vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13110__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16736_ clknet_leaf_140_wb_clk_i _02405_ _00965_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[709\]
+ sky130_fd_sc_hd__dfrtp_1
X_13948_ net1 team_04_WB.instance_to_wrap.wb_manage.curr_state\[1\] team_04_WB.instance_to_wrap.wb_manage.curr_state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__or3b_1
XANTENNA__08955__S net897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13661__A1 net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12464__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_159_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13661__B2 _07691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16667_ clknet_leaf_99_wb_clk_i _02336_ _00896_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[640\]
+ sky130_fd_sc_hd__dfrtp_1
X_13879_ _02921_ _03261_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15618_ net1240 vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__inv_2
XANTENNA__12216__A2 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16598_ clknet_leaf_13_wb_clk_i _02267_ _00827_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[571\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10227__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15549_ net1153 vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[44\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[12\]
+ net873 vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_170_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _03608_ net752 vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13177__B1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17219_ net1425 _02829_ _01465_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12924__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[809\] vssd1 vssd1
+ vccd1 vccd1 net2139 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_170_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold713 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[607\] vssd1 vssd1
+ vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold724 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[342\] vssd1 vssd1
+ vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[481\] vssd1 vssd1
+ vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold746 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[668\] vssd1 vssd1
+ vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14126__C1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold757 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[602\] vssd1 vssd1
+ vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold768 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[826\] vssd1 vssd1
+ vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05581_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[139\] vssd1 vssd1
+ vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12940__S net320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[303\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[271\]
+ net964 vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout297_A _07683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[625\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[593\]
+ net896 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout1004_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08451__S0 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09026__S net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08785_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[434\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[402\]
+ net866 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17280__1336 vssd1 vssd1 vccd1 vccd1 _17280__1336/HI net1336 sky130_fd_sc_hd__conb_1
XFILLER_0_137_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout464_A _06203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13101__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15552__A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_140_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08718__X _04329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12387__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10696__A net905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A _04838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_70 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout729_A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09406_ net724 _05010_ net714 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13404__A1 team_04_WB.MEM_SIZE_REG_REG\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09337_ _03723_ _03782_ _03630_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o21ai_2
XANTENNA__13955__A2 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout517_X net517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09084__B2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_168_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1259_X net1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13800__A team_04_WB.ADDR_START_VAL_REG\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _04875_ _04876_ _04877_ _04878_ net786 net801 vssd1 vssd1 vccd1 vccd1 _04879_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_161_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13168__B1 net291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[765\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[733\]
+ net945 vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09199_ _04804_ _04809_ net722 vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__mux2_1
XANTENNA__08172__Y _03783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12915__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ net582 _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_75_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08105__S net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14117__C1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11161_ net286 _06644_ _06646_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_112_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10112_ team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[5\] _03724_ _04002_
+ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and3_1
XANTENNA__14132__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_164_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ net630 net628 net552 vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_164_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ _05549_ _05653_ net643 _03836_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__o2bb2a_1
X_14920_ net1117 vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08442__S0 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12694__A2 net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[8\] vssd1 vssd1 vccd1
+ vccd1 net1477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 team_04_WB.instance_to_wrap.final_design.VGA_data_control.ready_data\[18\]
+ vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 _02764_ vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A DAT_I[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ net1170 vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__inv_2
Xhold73 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[25\] vssd1 vssd1
+ vccd1 vccd1 net1510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[2\] vssd1
+ vssd1 vccd1 vccd1 net1521 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 net158 vssd1 vssd1 vccd1 vccd1 net1532 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _03179_ _03180_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__or3_1
XANTENNA__08775__S _03640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__B1 _03621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14782_ net1218 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__inv_2
X_11994_ net2567 net516 _07450_ net448 vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__a22o_1
XANTENNA__08114__A3 _03635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ clknet_leaf_100_wb_clk_i _02190_ _00750_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[494\]
+ sky130_fd_sc_hd__dfrtp_1
X_13733_ _07772_ _07804_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__xnor2_1
X_10945_ net630 _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__nor2_1
XANTENNA__08110__A1_N net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_4_5__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16452_ clknet_leaf_168_wb_clk_i _02121_ _00681_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[425\]
+ sky130_fd_sc_hd__dfrtp_1
X_13664_ _03046_ _03053_ team_04_WB.ADDR_START_VAL_REG\[3\] vssd1 vssd1 vccd1 vccd1
+ _03055_ sky130_fd_sc_hd__a21oi_1
X_10876_ _04643_ _06358_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15403_ net1120 vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__inv_2
XFILLER_0_144_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12615_ _07584_ net487 net414 net2213 vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ clknet_leaf_155_wb_clk_i _02052_ _00612_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[356\]
+ sky130_fd_sc_hd__dfrtp_1
X_13595_ _03498_ _05925_ net1102 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11957__A1 _07398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15334_ net1110 vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12546_ net2479 net261 net422 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11421__A3 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13159__B1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15265_ net1167 vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ net2263 net430 _07651_ net524 vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_4 _07402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12906__B1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_111_wb_clk_i _02673_ _01233_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[977\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11230__A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ team_04_WB.instance_to_wrap.final_design.VGA_data_control.VGA_request_address\[1\]
+ _03416_ _03364_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o21ai_1
X_11428_ _06505_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15196_ net1148 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__inv_2
XANTENNA__12045__B net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14108__C1 net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[0\] team_04_WB.instance_to_wrap.final_design.vga.h_current_state\[1\]
+ _03366_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__and3_1
X_11359_ net582 _06847_ net288 vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14541__A net1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__A2 net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08681__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14123__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__B net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ net1488 _06102_ net1032 vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__mux2_1
X_13029_ _07490_ net374 net307 net1694 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a22o_1
Xfanout1060 net1061 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__buf_2
XFILLER_0_174_36 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__buf_2
Xfanout1082 net1083 vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_2
Xfanout1093 team_04_WB.instance_to_wrap.final_design.reqhand.current_client\[2\] vssd1
+ vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_174_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08570_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[886\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[854\]
+ net851 vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
XANTENNA__08685__S net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ clknet_leaf_189_wb_clk_i _02388_ _00948_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[692\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11948__A1 team_04_WB.instance_to_wrap.CPU_DAT_O\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09122_ _04729_ _04730_ _04731_ _04732_ net837 net748 vssd1 vssd1 vccd1 vccd1 _04733_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13620__A _07039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09161__S1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[748\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[716\]
+ net921 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A _07258_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08004_ _03591_ _03599_ _03609_ _03612_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_114_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold510 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[50\] vssd1 vssd1
+ vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold521 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[583\] vssd1 vssd1
+ vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold532 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[337\] vssd1 vssd1
+ vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13570__B1 net1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold543 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[92\] vssd1 vssd1
+ vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[357\] vssd1 vssd1
+ vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12670__S net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold565 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[478\] vssd1 vssd1
+ vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1121_A net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[555\] vssd1 vssd1
+ vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 team_04_WB.instance_to_wrap.final_design.VGA_data_control.data_to_VGA\[20\]
+ vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__A2 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[885\] vssd1 vssd1
+ vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A _07482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08906_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[880\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[848\]
+ net863 vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__mux2_1
X_09886_ net661 _04526_ _04527_ net636 vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__o211ai_1
Xhold1210 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[30\] vssd1 vssd1
+ vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 team_04_WB.instance_to_wrap.final_design.VGA_adr\[1\] vssd1 vssd1 vccd1
+ vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08837_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[465\] _03656_ _04447_
+ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout846_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[562\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[530\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11636__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__A3 net469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08699_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[179\] team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[147\]
+ net935 vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
X_10730_ net632 net630 net552 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__mux2_1
XANTENNA__13928__A2 net1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ team_04_WB.instance_to_wrap.final_design.reqhand.instruction\[20\] net1016
+ net1012 team_04_WB.instance_to_wrap.CPU_DAT_O\[20\] vssd1 vssd1 vccd1 vccd1 _02748_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14626__A net1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_157_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14050__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[13\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11939__B2 _07403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ net656 net605 net218 vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__and3_1
X_13380_ team_04_WB.instance_to_wrap.final_design.VGA_adr\[8\] team_04_WB.MEM_SIZE_REG_REG\[10\]
+ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12061__B1 _07485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ _06133_ net1519 net1022 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__mux2_1
XANTENNA__12600__A2 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ net255 net671 vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and2_2
XFILLER_0_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11688__C _06257_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_163_wb_clk_i clknet_4_9__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_163_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_15050_ net1116 vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__inv_2
X_12262_ net256 net675 vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__and2_1
XFILLER_0_142_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11213_ net558 _06600_ _06601_ _06690_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__o31a_1
X_14001_ _05445_ _03308_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__or2_2
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ net258 net650 vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__and2_1
XANTENNA__14361__A net1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14105__A2 _07703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ net554 _06213_ _06241_ _06247_ _06631_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__o32a_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15952_ net1406 _01628_ _00179_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11075_ _03892_ net544 _06563_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08415__S0 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14030__A_N team_04_WB.instance_to_wrap.BUSY_O vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ _05577_ _05636_ _05575_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__o21a_1
X_14903_ net1226 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__inv_2
XFILLER_0_170_9 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10678__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_output131_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ clknet_leaf_98_wb_clk_i _01560_ _00110_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__dfrtp_1
X_14834_ net1244 vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13616__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12419__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14765_ net1210 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__inv_2
X_11977_ team_04_WB.instance_to_wrap.final_design.reqhand.data_from_UART\[1\] team_04_WB.instance_to_wrap.CPU_DAT_O\[1\]
+ net266 vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__mux2_1
XANTENNA__13092__A2 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ clknet_leaf_150_wb_clk_i _02173_ _00733_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[477\]
+ sky130_fd_sc_hd__dfrtp_1
X_13716_ team_04_WB.ADDR_START_VAL_REG\[11\] _03099_ _03103_ _03106_ vssd1 vssd1 vccd1
+ vccd1 _03107_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ _06403_ _06416_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__nand2b_1
X_14696_ net1117 vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16435_ clknet_leaf_188_wb_clk_i _02104_ _00664_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[408\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13647_ net1098 _03034_ net1045 team_04_WB.instance_to_wrap.final_design.CPU_instr_adr\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o2bb2a_1
X_10859_ _04218_ _06347_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_1
XANTENNA__14536__A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14041__B2 team_04_WB.instance_to_wrap.CPU_DAT_O\[22\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16366_ clknet_leaf_27_wb_clk_i _02035_ _00595_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[339\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13578_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10783__B _06207_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15317_ net1207 vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__inv_2
X_12529_ net2363 net241 net420 vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__mux2_1
X_16297_ clknet_leaf_102_wb_clk_i _01966_ _00526_ vssd1 vssd1 vccd1 vccd1 team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[270\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15248_ net1163 vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10366__B1 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ net1128 vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09365__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_4
Xfanout319 _07675_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__B2 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ team_04_WB.instance_to_wrap.final_design.cpu.reg_window\[480\] _03650_ _03652_
+ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__or3_1
.ends

