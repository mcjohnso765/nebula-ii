* NGSPICE file created from team_10_Wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt team_10_Wrapper ACK_I ADR_O[0] ADR_O[10] ADR_O[11] ADR_O[12] ADR_O[13] ADR_O[14]
+ ADR_O[15] ADR_O[16] ADR_O[17] ADR_O[18] ADR_O[19] ADR_O[1] ADR_O[20] ADR_O[21] ADR_O[22]
+ ADR_O[23] ADR_O[24] ADR_O[25] ADR_O[26] ADR_O[27] ADR_O[28] ADR_O[29] ADR_O[2] ADR_O[30]
+ ADR_O[31] ADR_O[3] ADR_O[4] ADR_O[5] ADR_O[6] ADR_O[7] ADR_O[8] ADR_O[9] CYC_O DAT_I[0]
+ DAT_I[10] DAT_I[11] DAT_I[12] DAT_I[13] DAT_I[14] DAT_I[15] DAT_I[16] DAT_I[17]
+ DAT_I[18] DAT_I[19] DAT_I[1] DAT_I[20] DAT_I[21] DAT_I[22] DAT_I[23] DAT_I[24] DAT_I[25]
+ DAT_I[26] DAT_I[27] DAT_I[28] DAT_I[29] DAT_I[2] DAT_I[30] DAT_I[31] DAT_I[3] DAT_I[4]
+ DAT_I[5] DAT_I[6] DAT_I[7] DAT_I[8] DAT_I[9] DAT_O[0] DAT_O[10] DAT_O[11] DAT_O[12]
+ DAT_O[13] DAT_O[14] DAT_O[15] DAT_O[16] DAT_O[17] DAT_O[18] DAT_O[19] DAT_O[1] DAT_O[20]
+ DAT_O[21] DAT_O[22] DAT_O[23] DAT_O[24] DAT_O[25] DAT_O[26] DAT_O[27] DAT_O[28]
+ DAT_O[29] DAT_O[2] DAT_O[30] DAT_O[31] DAT_O[3] DAT_O[4] DAT_O[5] DAT_O[6] DAT_O[7]
+ DAT_O[8] DAT_O[9] SEL_O[0] SEL_O[1] SEL_O[2] SEL_O[3] STB_O WE_O gpio_in[0] gpio_in[10]
+ gpio_in[11] gpio_in[12] gpio_in[13] gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17]
+ gpio_in[18] gpio_in[19] gpio_in[1] gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23]
+ gpio_in[24] gpio_in[25] gpio_in[26] gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2]
+ gpio_in[30] gpio_in[31] gpio_in[32] gpio_in[33] gpio_in[34] gpio_in[35] gpio_in[36]
+ gpio_in[37] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[34]
+ gpio_oeb[35] gpio_oeb[36] gpio_oeb[37] gpio_oeb[3] gpio_oeb[4] gpio_oeb[5] gpio_oeb[6]
+ gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0] gpio_out[10] gpio_out[11] gpio_out[12]
+ gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16] gpio_out[17] gpio_out[18] gpio_out[19]
+ gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22] gpio_out[23] gpio_out[24] gpio_out[25]
+ gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29] gpio_out[2] gpio_out[30] gpio_out[31]
+ gpio_out[32] gpio_out[33] gpio_out[34] gpio_out[35] gpio_out[36] gpio_out[37] gpio_out[3]
+ gpio_out[4] gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] irq[0] irq[1]
+ irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[3] la_data_in[4] la_data_in[5] la_data_in[6]
+ la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10] la_data_out[11]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[3] la_data_out[4] la_data_out[5] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[3] la_oenb[4]
+ la_oenb[5] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__2479__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155_ _1564_ _1583_ _0906_ _1562_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_38_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2106_ team_10_WB.instance_to_wrap.dispFSM.guesses\[6\] net112 net138 net671 vssd1
+ vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3086_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _1537_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[79\] sky130_fd_sc_hd__mux2_1
X_2037_ team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] net110 net137 team_10_WB.instance_to_wrap.dispFSM.msg\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__o22a_1
XANTENNA__3050__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3443__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4670__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3988_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[25\]
+ _0056_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2939_ net214 net151 net120 net655 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[44\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_44_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2954__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2190__A team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout215_X net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4609_ net384 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_60_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4108__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4258__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4580__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1996__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3924__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2275__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3425__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3911_ net278 vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1987__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3842_ net242 vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2936__A1 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3773_ net272 vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2724_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ _1351_ team_10_WB.instance_to_wrap.clock_div.count\[9\] vssd1 vssd1 vccd1 vccd1
+ _1355_ sky130_fd_sc_hd__a31o_1
XANTENNA__3393__X _1770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2655_ _1308_ _1310_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4325_ clknet_leaf_14_wb_clk_i _0715_ _0314_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[48\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2586_ _0888_ _0902_ vssd1 vssd1 vccd1 vccd1 _1271_ sky130_fd_sc_hd__nand2_1
XANTENNA__4400__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout138 net142 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_2
X_4256_ clknet_leaf_0_wb_clk_i _0650_ _0245_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.green
+ sky130_fd_sc_hd__dfrtp_1
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_4
X_4187_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[49\]
+ _0176_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[49\] sky130_fd_sc_hd__dfrtp_1
X_3207_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] _1621_ vssd1 vssd1 vccd1
+ vccd1 _1622_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3138_ _1549_ _1567_ _1568_ _1551_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1
+ vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__o32a_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3416__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__mux2_1
XANTENNA__4173__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1978__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3744__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\] vssd1 vssd1 vccd1 vccd1
+ net627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 team_10_WB.instance_to_wrap.dispFSM.guesses\[64\] vssd1 vssd1 vccd1 vccd1
+ net638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2794__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3407__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3919__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1969__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4423__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ net545 net133 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\]
+ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3343__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2371_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] _1084_ _1144_
+ _1145_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__o22a_1
X_4110_ clknet_leaf_18_wb_clk_i net500 _0109_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_4041_ clknet_leaf_19_wb_clk_i _0526_ _0082_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1902__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_1054 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3829__A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3825_ net256 vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__inv_2
XANTENNA__2452__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3756_ net286 vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__inv_2
X_2707_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1 _1345_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3687_ net244 vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3564__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2638_ _0922_ _0925_ _0935_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] _0975_
+ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__o221a_1
XANTENNA__2252__A_N team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2569_ net223 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] net227 vssd1
+ vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__and3_1
X_4308_ clknet_leaf_18_wb_clk_i net574 _0297_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4239_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[3\]
+ _0228_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__4168__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4446__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1940_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] net147 vssd1 vssd1 vccd1
+ vccd1 _0863_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1871_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] vssd1 vssd1 vccd1 vccd1
+ _0796_ sky130_fd_sc_hd__inv_2
X_4590_ net454 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
X_3610_ net263 vssd1 vssd1 vccd1 vccd1 _0142_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3541_ net236 vssd1 vssd1 vccd1 vccd1 _0073_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3472_ team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] _1715_ _1842_ _0821_ vssd1
+ vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__a211o_1
X_2423_ net469 net129 vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__or2_1
XANTENNA__3963__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2354_ _1126_ _1128_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2285_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _1063_ _1064_ _1066_ vssd1
+ vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__a22o_1
XANTENNA__2447__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4024_ clknet_leaf_0_wb_clk_i net473 _0071_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4469__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3808_ net293 vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_586 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3739_ net272 vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__inv_2
X_4690__438 vssd1 vssd1 vccd1 vccd1 _4690__438/HI net438 sky130_fd_sc_hd__conb_1
XFILLER_0_28_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input2_X net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3188__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3932__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2070_ team_10_WB.instance_to_wrap.dispFSM.guesses\[42\] net113 net140 net668 vssd1
+ vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_6_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3482__B1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] _0835_ net160 vssd1 vssd1 vccd1
+ vccd1 _1487_ sky130_fd_sc_hd__a41o_1
XFILLER_0_56_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1923_ net4 net5 net300 vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__o21ba_1
X_4642_ net411 vssd1 vssd1 vccd1 vccd1 la_data_out[12] sky130_fd_sc_hd__buf_2
XANTENNA__4271__Q team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ net449 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3524_ net245 vssd1 vssd1 vccd1 vccd1 _0056_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3455_ team_10_WB.instance_to_wrap.host_row2\[54\] net170 net167 team_10_WB.instance_to_wrap.host_row2\[78\]
+ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload27_A clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4141__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2406_ team_10_WB.instance_to_wrap.clock_div.count\[19\] team_10_WB.instance_to_wrap.clock_div.count\[18\]
+ team_10_WB.instance_to_wrap.clock_div.count\[21\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__or4_1
X_3386_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1704_ net179 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\]
+ _1762_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout192_A _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2337_ _0809_ _0866_ _1093_ _0811_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__a22oi_1
XANTENNA__3053__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2268_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0800_ net215 _0792_ vssd1
+ vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_4_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4673__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4291__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ clknet_leaf_23_wb_clk_i _0495_ net274 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_2199_ _0984_ _0987_ _0975_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_36_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2640__B net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2200__A1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3752__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold41 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] vssd1 vssd1 vccd1 vccd1
+ net498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 team_10_WB.instance_to_wrap.gamelogic.red vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 team_10_WB.instance_to_wrap.host_row1\[72\] vssd1 vssd1 vccd1 vccd1 net531
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 net520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold52 _0674_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 team_10_WB.instance_to_wrap.host_row1\[41\] vssd1 vssd1 vccd1 vccd1 net553
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] vssd1 vssd1 vccd1
+ vccd1 net542 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input18_A wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3464__B1 _1837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4014__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_35_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_5 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4164__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3240_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\] _1642_ net172 vssd1
+ vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__a21oi_1
X_3171_ _1550_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__nor2_1
X_2122_ net219 net218 team_10_WB.instance_to_wrap.gamelogic.state\[2\] team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__or4b_2
XANTENNA__3455__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2258__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2053_ team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] net110 net137 net605 vssd1
+ vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2955_ _0798_ _1478_ net159 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[7\] sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1906_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _0829_ sky130_fd_sc_hd__inv_2
X_2886_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] net1 _1467_ vssd1 vssd1 vccd1
+ vccd1 _1468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4625_ team_10_WB.instance_to_wrap.lcdPlayer.lcd_en vssd1 vssd1 vccd1 vccd1 net77
+ sky130_fd_sc_hd__clkbuf_1
X_4556_ net368 vssd1 vssd1 vccd1 vccd1 DAT_O[30] sky130_fd_sc_hd__buf_2
XANTENNA_fanout205_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2194__B1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3507_ net246 vssd1 vssd1 vccd1 vccd1 _0039_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4668__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4487_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[44\]
+ _0470_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_12_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3438_ _1719_ _1801_ _1810_ net179 vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ team_10_WB.instance_to_wrap.host_row1\[50\] _1699_ net167 team_10_WB.instance_to_wrap.host_row2\[74\]
+ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__a22o_1
XANTENNA__2249__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3446__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4037__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4187__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3382__C1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[12] sky130_fd_sc_hd__buf_2
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_0_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1999__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2740_ team_10_WB.instance_to_wrap.clock_div.count\[13\] team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ team_10_WB.instance_to_wrap.clock_div.count\[15\] _1362_ vssd1 vssd1 vccd1 vccd1
+ _1365_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2671_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] _1324_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[7\]
+ _0393_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4341_ clknet_leaf_16_wb_clk_i _0731_ _0330_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[64\]
+ sky130_fd_sc_hd__dfstp_1
X_4272_ clknet_leaf_0_wb_clk_i _0662_ _0261_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3223_ net172 _1631_ _1632_ vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__nor3_1
XFILLER_0_20_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3154_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] _0899_ _1582_ vssd1
+ vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_38_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3428__B1 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2105_ team_10_WB.instance_to_wrap.dispFSM.guesses\[15\] net145 _0915_ net508 vssd1
+ vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__a22o_1
X_3085_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__mux2_1
X_2036_ team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] net113 net141 team_10_WB.instance_to_wrap.dispFSM.msg\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0743_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout155_A _1182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3987_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[24\]
+ _0055_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3567__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2938_ net215 net151 net120 net664 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[43\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4502__314 vssd1 vssd1 vccd1 vccd1 _4502__314/HI net314 sky130_fd_sc_hd__conb_1
XANTENNA__2190__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2869_ team_10_WB.instance_to_wrap.host_message_reg.Cstate net157 _1302_ vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.next_state sky130_fd_sc_hd__a21o_1
X_4608_ net383 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_fanout208_X net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4539_ net351 vssd1 vssd1 vccd1 vccd1 DAT_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_7_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_392 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3355__C1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3370__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4202__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3940__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4352__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3910_ net259 vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3841_ net241 vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2291__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3772_ net291 vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__inv_2
XANTENNA__2936__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2723_ net731 _1354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[8\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2654_ _1228_ _1309_ _1315_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
X_2585_ _1265_ _1269_ vssd1 vssd1 vccd1 vccd1 _1270_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3361__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4324_ clknet_leaf_18_wb_clk_i net559 _0313_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout117 net119 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_2
Xfanout128 _1188_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4255_ clknet_leaf_14_wb_clk_i _0649_ _0244_ vssd1 vssd1 vccd1 vccd1 team_10_WB.EN_VAL_REG
+ sky130_fd_sc_hd__dfrtp_1
Xfanout139 net142 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__dlymetal6s2s_1
X_4186_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[48\]
+ _0175_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[48\] sky130_fd_sc_hd__dfrtp_1
X_3206_ _1621_ _1611_ _1620_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__and3b_1
XANTENNA__3061__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137_ _1275_ _1550_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__or2_1
X_4647__416 vssd1 vssd1 vccd1 vccd1 _4647__416/HI net416 sky130_fd_sc_hd__conb_1
X_3068_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] _1528_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[70\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2019_ _0890_ net228 net222 vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2388__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4225__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3352__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[13\] vssd1 vssd1
+ vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _0722_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] vssd1 vssd1 vccd1 vccd1
+ net650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] vssd1 vssd1 vccd1 vccd1
+ net639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4375__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4364__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2918__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3343__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1145_ sky130_fd_sc_hd__a21o_1
XANTENNA__3670__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ clknet_leaf_21_wb_clk_i _0525_ _0081_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4274__Q team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3824_ net248 vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__inv_2
XANTENNA__2909__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3755_ net272 vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2706_ net580 net546 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[1\]
+ sky130_fd_sc_hd__xor2_1
X_3686_ net234 vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2637_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _1085_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ _1303_ vssd1 vssd1 vccd1 vccd1 _0005_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout118_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2568_ _0974_ _1253_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4676__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2499_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] _1218_ _1217_ vssd1
+ vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__mux2_1
X_4307_ clknet_leaf_20_wb_clk_i _0697_ _0296_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_4238_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[2\]
+ _0227_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3098__A1 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4169_ clknet_leaf_26_wb_clk_i _0638_ _0158_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\]
+ sky130_fd_sc_hd__dfstp_2
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4508__320 vssd1 vssd1 vccd1 vccd1 _4508__320/HI net320 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_61_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3325__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1870_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] vssd1 vssd1 vccd1 vccd1
+ _0795_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3665__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3540_ net236 vssd1 vssd1 vccd1 vccd1 _0072_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3471_ team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] net173 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[15\]
+ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a221o_1
X_2422_ net158 _1181_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2353_ _1099_ _1124_ _1125_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__or3_1
XANTENNA__4269__Q team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2284_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _1065_ vssd1 vssd1 vccd1
+ vccd1 _1066_ sky130_fd_sc_hd__xnor2_1
X_4023_ clknet_leaf_0_wb_clk_i net471 _0070_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4070__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout235_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ net281 vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1999_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] net148 net118
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] vssd1 vssd1 vccd1 vccd1 _0750_
+ sky130_fd_sc_hd__o22a_1
X_3738_ net295 vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3669_ net240 vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4413__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3467__D1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\] _0834_ net164 vssd1 vssd1 vccd1
+ vccd1 _1486_ sky130_fd_sc_hd__a41o_1
XFILLER_0_56_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1922_ net304 net5 vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4641_ net410 vssd1 vssd1 vccd1 vccd1 la_data_out[11] sky130_fd_sc_hd__buf_2
XFILLER_0_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4572_ net448 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XFILLER_0_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3523_ net245 vssd1 vssd1 vccd1 vccd1 _0055_ sky130_fd_sc_hd__inv_2
X_3454_ team_10_WB.instance_to_wrap.host_row1\[70\] _1703_ net179 team_10_WB.instance_to_wrap.host_row2\[70\]
+ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2405_ team_10_WB.instance_to_wrap.clock_div.count\[14\] team_10_WB.instance_to_wrap.clock_div.count\[17\]
+ team_10_WB.instance_to_wrap.clock_div.count\[16\] team_10_WB.instance_to_wrap.clock_div.count\[15\]
+ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3385_ team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] net171 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4436__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2336_ _1103_ _1104_ _1105_ _1106_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_4_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2458__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2267_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] _0801_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout185_A _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4006_ clknet_leaf_23_wb_clk_i _0494_ net274 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2276__A2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2198_ _0976_ _0977_ _0980_ _0985_ _0986_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2433__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold31 team_10_WB.instance_to_wrap.message_reg.msg\[0\] vssd1 vssd1 vccd1 vccd1 net488
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 _0506_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] vssd1 vssd1 vccd1 vccd1
+ net510 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 team_10_WB.instance_to_wrap.host_row1\[45\] vssd1 vssd1 vccd1 vccd1 net499
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 team_10_WB.instance_to_wrap.message_reg.msg\[1\] vssd1 vssd1 vccd1 vccd1 net521
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] vssd1 vssd1 vccd1
+ vccd1 net554 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 team_10_WB.instance_to_wrap.clock_div.count\[27\] vssd1 vssd1 vccd1 vccd1
+ net532 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 team_10_WB.instance_to_wrap.message_reg.msg\[7\] vssd1 vssd1 vccd1 vccd1 net543
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4372__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3419__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4309__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3943__A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4459__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3170_ _0903_ _1277_ net195 vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__and3b_1
X_2121_ team_10_WB.instance_to_wrap.gamelogic.state\[2\] _0923_ team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__and3b_1
X_2052_ team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] net115 net135 net703 vssd1
+ vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_24_wb_clk_i_X clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2954_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\] net165 _1478_ net213 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[6\] sky130_fd_sc_hd__o22a_1
X_1905_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0828_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2885_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] vssd1 vssd1 vccd1 vccd1
+ _1467_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4624_ net394 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4555_ net367 vssd1 vssd1 vccd1 vccd1 DAT_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_12_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3391__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3506_ net245 vssd1 vssd1 vccd1 vccd1 _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4486_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[43\]
+ _0469_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3437_ _1799_ _1803_ _1808_ _1811_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__or4_1
X_3368_ net610 net177 _1746_ net230 vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_51_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2188__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4684__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2319_ _0867_ _1090_ vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__or2_1
X_3299_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__or2_1
XANTENNA__3976__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3382__B1 _1752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2488__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[13] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_17 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1999__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2948__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4131__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2670_ _1324_ _1325_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4281__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3373__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1923__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4340_ clknet_leaf_19_wb_clk_i _0730_ _0329_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_4271_ clknet_leaf_0_wb_clk_i _0661_ _0260_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3222_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ _1628_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2479__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3153_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\]
+ net228 vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o21a_1
XANTENNA__3999__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2104_ team_10_WB.instance_to_wrap.dispFSM.guesses\[8\] net114 net141 net695 vssd1
+ vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4569__445 vssd1 vssd1 vccd1 vccd1 net445 _4569__445/LO sky130_fd_sc_hd__conb_1
X_3084_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] _1536_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[78\] sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4005__RESET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2035_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] net143 net107 net678 vssd1 vssd1
+ vccd1 vccd1 _0744_ sky130_fd_sc_hd__a22o_1
XANTENNA__3848__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2939__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3986_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[23\]
+ _0054_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout148_A net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2937_ net216 net151 net120 net677 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[42\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3059__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4541__353 vssd1 vssd1 vccd1 vccd1 _4541__353/HI net353 sky130_fd_sc_hd__conb_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4607_ net382 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2868_ net506 _1455_ _1440_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__4679__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2799_ _1407_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4538_ net350 vssd1 vssd1 vccd1 vccd1 DAT_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[26\]
+ _0452_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4154__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4525__337 vssd1 vssd1 vccd1 vccd1 _4525__337/HI net337 sky130_fd_sc_hd__conb_1
XFILLER_0_55_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3310__D_N net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ net241 vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3771_ net271 vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2722_ _1180_ _1353_ _1354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2653_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] _0827_ _1225_ _1233_
+ _1313_ vssd1 vssd1 vccd1 vccd1 _1315_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3346__B1 _1713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2584_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4027__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4323_ clknet_leaf_20_wb_clk_i _0713_ _0312_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout107 net108 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
Xfanout129 _1184_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
X_4254_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[10\]
+ _0243_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3205_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] _1392_ vssd1 vssd1 vccd1 vccd1
+ _1621_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4177__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4185_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[47\]
+ _0174_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[47\] sky130_fd_sc_hd__dfrtp_1
X_4612__387 vssd1 vssd1 vccd1 vccd1 _4612__387/HI net387 sky130_fd_sc_hd__conb_1
X_3136_ _0903_ _1566_ _1280_ _1277_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__o211a_1
X_3067_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1528_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout265_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _0892_ net232 net2 vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_46_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3969_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[6\]
+ _0037_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold161 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\] vssd1 vssd1 vccd1 vccd1
+ net618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold150 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] vssd1 vssd1 vccd1 vccd1
+ net607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1
+ net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\] vssd1 vssd1 vccd1
+ vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] vssd1 vssd1 vccd1 vccd1
+ net640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4380__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3427__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2000__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3823_ net258 vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__inv_2
XANTENNA__3016__C1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3754_ net282 vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_9_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3685_ net244 vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_279 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2705_ net546 _1171_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2636_ net160 _1301_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2567_ _1047_ _1252_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1
+ vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2498_ _0812_ _0888_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__nor2_1
X_4306_ clknet_leaf_19_wb_clk_i _0696_ _0295_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3072__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4237_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[1\]
+ _0226_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] sky130_fd_sc_hd__dfrtp_1
X_4168_ clknet_leaf_25_wb_clk_i _0637_ _0157_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4099_ clknet_leaf_12_wb_clk_i _0570_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout170_X net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1278_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__and3b_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3022__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4342__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4492__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4199__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3470_ team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] net175 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__a22o_1
X_2421_ net162 net154 vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__nor2_1
X_2352_ _1117_ _1122_ _1127_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__and3_1
XANTENNA__2524__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2283_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__nand2_1
X_4022_ clknet_leaf_0_wb_clk_i net482 _0069_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4683__436 vssd1 vssd1 vccd1 vccd1 _4683__436/HI net436 sky130_fd_sc_hd__conb_1
XANTENNA__4215__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_414 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout130_A net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3806_ net294 vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4365__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3737_ net292 vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1998_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] net148 net118
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1 _0751_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_697 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3668_ net277 vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__inv_2
XANTENNA__4687__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3599_ net276 vssd1 vssd1 vccd1 vccd1 _0131_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2619_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_54_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2451__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_14_wb_clk_i_X clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout290 net291 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__buf_4
XANTENNA_clkload6_A clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4388__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _0835_ net160 vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1921_ net300 net4 vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__and2b_1
XANTENNA__2442__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ net409 vssd1 vssd1 vccd1 vccd1 la_data_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_56_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2993__B2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4571_ net447 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3522_ net245 vssd1 vssd1 vccd1 vccd1 _0054_ sky130_fd_sc_hd__inv_2
X_3453_ team_10_WB.instance_to_wrap.host_row2\[86\] _1686_ _1695_ net302 vssd1 vssd1
+ vccd1 vccd1 _1827_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_667 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2404_ _1165_ _1166_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3384_ net66 net178 _1761_ net230 vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2335_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\] _1089_ vssd1 vssd1
+ vccd1 vccd1 _1111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2266_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] net217 vssd1 vssd1 vccd1
+ vccd1 _1048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4005_ clknet_leaf_23_wb_clk_i _0493_ net274 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2197_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] net212 vssd1 vssd1 vccd1
+ vccd1 _0986_ sky130_fd_sc_hd__xor2_1
XANTENNA__3473__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2433__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3161__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold32 team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net489
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\] vssd1 vssd1 vccd1 vccd1
+ net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] vssd1 vssd1 vccd1 vccd1 net467
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _0581_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 team_10_WB.instance_to_wrap.host_row1\[79\] vssd1 vssd1 vccd1 vccd1 net511
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] vssd1 vssd1 vccd1
+ vccd1 net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 team_10_WB.instance_to_wrap.host_row1\[52\] vssd1 vssd1 vccd1 vccd1 net544
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 team_10_WB.instance_to_wrap.host_row1\[59\] vssd1 vssd1 vccd1 vccd1 net555
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net533 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_51_Left_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3496__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2975__B2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_7 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_829 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3435__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4060__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2120_ net219 net218 vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_23_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2051_ team_10_WB.instance_to_wrap.dispFSM.guesses\[69\] net143 net107 net569 vssd1
+ vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__a22o_1
XANTENNA__3455__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1134 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2953_ _0800_ _1478_ _1474_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[5\]
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_33_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1904_ net242 vssd1 vssd1 vccd1 vccd1 _0018_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2884_ net193 _1466_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[4\]
+ sky130_fd_sc_hd__and2_1
X_4623_ team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs vssd1 vssd1 vccd1 vccd1 net76
+ sky130_fd_sc_hd__buf_1
XFILLER_0_4_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4554_ net366 vssd1 vssd1 vccd1 vccd1 DAT_O[28] sky130_fd_sc_hd__buf_2
XFILLER_0_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4403__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3391__A1 team_10_WB.instance_to_wrap.host_row2\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3505_ net250 vssd1 vssd1 vccd1 vccd1 _0037_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4485_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[42\]
+ _0468_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3436_ _1715_ _1720_ _0821_ team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1
+ vccd1 vccd1 _1811_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ net179 _1744_ _1745_ _1743_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_51_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2318_ team_10_WB.instance_to_wrap.host_col\[3\] _0868_ _1092_ _0846_ _0856_ vssd1
+ vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__o311ai_1
X_3298_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__nor2_1
XANTENNA__3080__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2249_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] _0799_ net214 _0794_ _1030_
+ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__a221o_1
XANTENNA__3446__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3382__B2 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__clkbuf_4
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput44 net44 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[15] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_737 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2948__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4426__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1923__A2 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4270_ clknet_leaf_0_wb_clk_i _0660_ _0259_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3221_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ net718 vssd1
+ vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__a21oi_1
X_3152_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] _1290_ _1550_ _1283_ vssd1 vssd1
+ vccd1 vccd1 _1581_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2103_ team_10_WB.instance_to_wrap.dispFSM.guesses\[9\] net110 net137 net662 vssd1
+ vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__o22a_1
XANTENNA__1921__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3083_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3428__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2034_ team_10_WB.instance_to_wrap.dispFSM.guesses\[78\] net112 net138 team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2939__A1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3985_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[22\]
+ _0053_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2936_ net217 net155 net123 net652 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[41\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_44_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2867_ _1455_ _1456_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[9\]
+ sky130_fd_sc_hd__nor2_1
X_4606_ net381 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2798_ _0815_ net177 _1406_ net282 vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__a211o_2
X_4537_ net349 vssd1 vssd1 vccd1 vccd1 DAT_O[11] sky130_fd_sc_hd__buf_2
XANTENNA__3075__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4468_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[25\]
+ _0451_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
X_3419_ team_10_WB.instance_to_wrap.host_row2\[68\] team_10_WB.instance_to_wrap.dispFSM.guesses\[44\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__mux2_1
XANTENNA__3116__A1 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4399_ clknet_leaf_5_wb_clk_i _0784_ _0382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_36_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2943__A team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3052__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3770_ net295 vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2721_ team_10_WB.instance_to_wrap.clock_div.count\[7\] _1351_ vssd1 vssd1 vccd1
+ vccd1 _1354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2652_ _1313_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2583_ _1256_ _1258_ _1266_ _1267_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3966__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4322_ clknet_leaf_25_wb_clk_i net566 _0311_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout119 _0875_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_2
X_4253_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[9\]
+ _0242_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout108 _0915_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
X_3204_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\] _1619_ vssd1 vssd1 vccd1
+ vccd1 _1620_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4184_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[46\]
+ _0173_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[46\] sky130_fd_sc_hd__dfrtp_1
X_3135_ _1561_ _1565_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__xnor2_1
X_3066_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _1527_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\] sky130_fd_sc_hd__mux2_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2017_ net2 net301 _0893_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2482__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3968_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[5\]
+ _0036_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3034__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2919_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\] net152 net120 net722
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[24\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3899_ net254 vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout213_X net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\] vssd1 vssd1 vccd1
+ vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\] vssd1 vssd1 vccd1
+ vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] vssd1 vssd1 vccd1 vccd1
+ net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 net69 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] vssd1 vssd1 vccd1
+ vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] vssd1 vssd1 vccd1 vccd1
+ net641 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4121__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3025__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3009__A team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2000__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3822_ net258 vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3753_ net292 vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2704_ team_10_WB.instance_to_wrap.host_col\[3\] net220 net300 vssd1 vssd1 vccd1
+ vccd1 net81 sky130_fd_sc_hd__mux2_1
X_3684_ net237 vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2635_ _0841_ _1086_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__nor2_2
XANTENNA__4144__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4653__422 vssd1 vssd1 vccd1 vccd1 _4653__422/HI net422 sky130_fd_sc_hd__conb_1
X_4305_ clknet_leaf_12_wb_clk_i _0695_ _0294_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_2566_ net218 _0948_ net134 vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__o21ai_1
X_2497_ net220 _0891_ _1217_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4294__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4236_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[0\]
+ _0225_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4167_ clknet_leaf_25_wb_clk_i _0636_ _0156_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3098__A3 _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3118_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] _1278_ vssd1 vssd1 vccd1 vccd1
+ _1549_ sky130_fd_sc_hd__and2_1
X_4098_ clknet_leaf_12_wb_clk_i _0569_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_3049_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1519_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3101__B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_18 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4017__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3011__B net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4167__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4637__406 vssd1 vssd1 vccd1 vccd1 _4637__406/HI net406 sky130_fd_sc_hd__conb_1
XFILLER_0_49_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1980__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2420_ net202 _0942_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2351_ _1094_ _1097_ net225 _0869_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__o2bb2a_1
X_2282_ _0990_ _1063_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nor2_1
X_4021_ clknet_leaf_0_wb_clk_i net477 _0068_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3348__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3805_ net287 vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__inv_2
X_1997_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] net148 net118
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] vssd1 vssd1 vccd1 vccd1 _0752_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3736_ net293 vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3667_ net259 vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3598_ net261 vssd1 vssd1 vccd1 vccd1 _0130_ sky130_fd_sc_hd__inv_2
X_2618_ _1294_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\] _1074_ vssd1 vssd1
+ vccd1 vccd1 _0006_ sky130_fd_sc_hd__mux2_1
X_2549_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\]
+ _1240_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\] vssd1 vssd1
+ vccd1 vccd1 _1241_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_54_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4219_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[81\]
+ _0208_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[81\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3476__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout280 net282 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_4
Xfanout291 net299 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1920_ net304 net2 vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4570_ net446 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XFILLER_0_4_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3521_ net245 vssd1 vssd1 vccd1 vccd1 _0053_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2800__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3452_ team_10_WB.instance_to_wrap.host_row1\[54\] _1699_ net180 team_10_WB.instance_to_wrap.host_row2\[62\]
+ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3383_ net303 _1758_ _1759_ net169 _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__a221o_1
X_2403_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ team_10_WB.instance_to_wrap.clock_div.count\[25\] team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2334_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\] _0868_ vssd1 vssd1
+ vccd1 vccd1 _1110_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2265_ _1035_ _1040_ _1046_ _0949_ vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__a31o_1
XANTENNA__3458__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2196_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _0801_ _0978_ _0979_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__a221o_1
X_4004_ clknet_leaf_23_wb_clk_i _0492_ net270 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2130__A0 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4332__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout240_A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4482__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3078__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout126_X net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3719_ net237 vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2011__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] vssd1 vssd1 vccd1 vccd1 net479
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 _0510_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\] vssd1 vssd1 vccd1 vccd1
+ net512 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\] vssd1 vssd1 vccd1
+ vccd1 net490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[7\] vssd1 vssd1 vccd1 vccd1
+ net501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__B1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 team_10_WB.instance_to_wrap.host_row1\[73\] vssd1 vssd1 vccd1 vccd1 net545
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold99 team_10_WB.instance_to_wrap.clock_div.count\[4\] vssd1 vssd1 vccd1 vccd1 net556
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[1\] vssd1 vssd1
+ vccd1 vccd1 net534 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 team_10_WB.instance_to_wrap.host_row1\[56\] vssd1 vssd1 vccd1 vccd1 net523
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4205__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4355__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] net111 net139 team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2952_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] net165 _1478_ net214 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[4\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_33_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3687__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2415__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1903_ team_10_WB.instance_to_wrap.uart_receiver.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2883_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] _1465_ vssd1 vssd1 vccd1
+ vccd1 _1466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4622_ team_10_WB.instance_to_wrap.uart_transmitter.tx_serial vssd1 vssd1 vccd1 vccd1
+ net75 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4553_ net365 vssd1 vssd1 vccd1 vccd1 DAT_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4484_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[41\]
+ _0467_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3391__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3504_ net251 vssd1 vssd1 vccd1 vccd1 _0036_ sky130_fd_sc_hd__inv_2
XANTENNA__2530__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3435_ team_10_WB.instance_to_wrap.host_row2\[69\] team_10_WB.instance_to_wrap.dispFSM.guesses\[45\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload25_A clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ net210 _0817_ _1690_ _1403_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_51_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ net510 _1677_ _1678_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout190_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2317_ net229 _0848_ _0855_ team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1
+ vccd1 vccd1 _1093_ sky130_fd_sc_hd__o211a_1
X_2248_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] _0801_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2103__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2179_ team_10_WB.instance_to_wrap.correct\[0\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__clkbuf_4
X_4592__456 vssd1 vssd1 vccd1 vccd1 net456 _4592__456/LO sky130_fd_sc_hd__conb_1
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput45 net45 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4378__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[16] sky130_fd_sc_hd__clkbuf_4
XANTENNA__2947__Y _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2203__X _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3373__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3220_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ _1630_ vssd1
+ vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3151_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] _1551_ _1579_ _1580_ vssd1 vssd1
+ vccd1 vccd1 _0497_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2102_ team_10_WB.instance_to_wrap.dispFSM.guesses\[10\] net114 net142 net694 vssd1
+ vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o22a_1
X_3082_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _1535_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[77\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2033_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] net144 net108 net595 vssd1 vssd1
+ vccd1 vccd1 _0746_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3984_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[21\]
+ _0052_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_2935_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] net152 net121 net696 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[40\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_44_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2866_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] _1454_ net176
+ vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__o21ai_1
X_4605_ net380 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_5_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2797_ team_10_WB.instance_to_wrap.lcdPlayer.currentState\[3\] net177 vssd1 vssd1
+ vccd1 vccd1 _1406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4536_ net348 vssd1 vssd1 vccd1 vccd1 DAT_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_41_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4467_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[24\]
+ _0450_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_3418_ _1790_ _1793_ net303 vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o21a_1
X_4398_ clknet_leaf_5_wb_clk_i _0783_ _0381_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[35\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_input8_A wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3349_ _1680_ _1718_ net179 _1728_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3104__B net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4050__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3355__A2 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2563__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2720_ team_10_WB.instance_to_wrap.clock_div.count\[7\] _1351_ vssd1 vssd1 vccd1
+ vccd1 _1353_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2651_ _1310_ _1312_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_10_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2582_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] _1259_ _0901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1267_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_10_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ clknet_leaf_10_wb_clk_i _0711_ _0310_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[44\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
X_4252_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[8\]
+ _0241_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3203_ _1619_ _1611_ _1618_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and3b_1
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4183_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[45\]
+ _0172_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[45\] sky130_fd_sc_hd__dfrtp_1
X_3134_ _1563_ _1564_ net221 _0906_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__o2bb2a_1
X_3065_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__mux2_1
XANTENNA__4073__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2016_ net4 _0887_ _0892_ net227 vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__or4b_2
XFILLER_0_49_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A _1182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3967_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[4\]
+ _0035_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2918_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\] net156 net125 net590
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[23\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__3875__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3898_ net258 vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2849_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\] _1442_ vssd1 vssd1
+ vccd1 vccd1 _1445_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout206_X net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_251 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4519_ net331 vssd1 vssd1 vccd1 vccd1 ADR_O[26] sky130_fd_sc_hd__buf_2
Xhold152 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\] vssd1 vssd1 vccd1
+ vccd1 net609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold130 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _0688_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1
+ net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1
+ net631 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\] vssd1 vssd1 vccd1
+ vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\] vssd1 vssd1 vccd1
+ vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4416__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531__343 vssd1 vssd1 vccd1 vccd1 _4531__343/HI net343 sky130_fd_sc_hd__conb_1
XANTENNA__4096__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3821_ net254 vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3695__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3752_ net299 vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3683_ net282 vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2703_ net225 net221 net300 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__mux2_1
XFILLER_0_40_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2634_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ _1083_ _1075_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__o31a_1
X_2565_ _0974_ _1251_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_40 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4304_ clknet_leaf_16_wb_clk_i _0694_ _0293_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4439__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2496_ net228 _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__nor2_1
X_4235_ clknet_leaf_21_wb_clk_i _0648_ _0224_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.state\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4166_ clknet_leaf_24_wb_clk_i _0635_ _0155_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3117_ net586 net5 _1548_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4097_ clknet_leaf_12_wb_clk_i _0568_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout270_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3048_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _1518_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[60\] sky130_fd_sc_hd__mux2_1
XFILLER_0_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout156_X net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_891 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4515__327 vssd1 vssd1 vccd1 vccd1 _4515__327/HI net327 sky130_fd_sc_hd__conb_1
XANTENNA__3956__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2049__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4602__377 vssd1 vssd1 vccd1 vccd1 _4602__377/HI net377 sky130_fd_sc_hd__conb_1
XFILLER_0_52_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__1980__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1980__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2350_ _1124_ _1125_ _1099_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__o21ai_1
X_2281_ _1012_ _1061_ _1062_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ clknet_leaf_0_wb_clk_i net480 _0067_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1002 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2460__A2 _1184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4111__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1996_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _0874_ _0884_ net158 vssd1
+ vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__o211a_1
XANTENNA__2533__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3804_ net287 vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3735_ net280 vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout116_A net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3666_ net271 vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3597_ net276 vssd1 vssd1 vccd1 vccd1 _0129_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2617_ _0830_ _1116_ _1119_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__nor3_1
X_2548_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_54_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4218_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[80\]
+ _0207_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[80\] sky130_fd_sc_hd__dfrtp_1
X_2479_ net544 net130 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__a22o_1
X_4149_ clknet_leaf_12_wb_clk_i _0620_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2451__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload0 clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2911__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3467__A1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_2
Xfanout292 net294 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 net274 vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_17_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4134__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2442__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4284__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3520_ net245 vssd1 vssd1 vccd1 vccd1 _0052_ sky130_fd_sc_hd__inv_2
X_3451_ net630 net177 _1825_ net230 vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3382_ net210 _1690_ _1752_ net232 _1403_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__a221o_1
X_2402_ team_10_WB.instance_to_wrap.clock_div.count\[27\] team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ team_10_WB.instance_to_wrap.clock_div.count\[29\] team_10_WB.instance_to_wrap.clock_div.count\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__or4_1
X_2333_ _0810_ _0843_ net196 vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2902__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2264_ _1038_ _1039_ _1041_ _1043_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__1940__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2195_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _0802_ _0981_ _0983_ vssd1
+ vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__o211a_1
X_4003_ clknet_leaf_24_wb_clk_i _0491_ net270 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_51 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2433__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1979_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net147 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout119_X net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3718_ net244 vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3649_ net264 vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold12 team_10_WB.instance_to_wrap.host_row1\[101\] vssd1 vssd1 vccd1 vccd1 net469
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2011__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 _0505_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _0547_ vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[1\] vssd1 vssd1
+ vccd1 vccd1 net491 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold45 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[7\] vssd1 vssd1 vccd1
+ vccd1 net502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 team_10_WB.instance_to_wrap.host_row1\[50\] vssd1 vssd1 vccd1 vccd1 net535
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold89 team_10_WB.instance_to_wrap.clock_div.count\[0\] vssd1 vssd1 vccd1 vccd1 net546
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4157__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 team_10_WB.instance_to_wrap.message_reg.msg\[6\] vssd1 vssd1 vccd1 vccd1 net524
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3385__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2951_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] net162 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[3\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_33_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4608__383 vssd1 vssd1 vccd1 vccd1 _4608__383/HI net383 sky130_fd_sc_hd__conb_1
XFILLER_0_32_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1902_ net202 vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__inv_2
X_4621_ net393 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XFILLER_0_38_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2882_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net224 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__or3b_1
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3376__B1 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4552_ net364 vssd1 vssd1 vccd1 vccd1 DAT_O[26] sky130_fd_sc_hd__buf_2
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4483_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[40\]
+ _0466_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3503_ net250 vssd1 vssd1 vccd1 vccd1 _0035_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3434_ team_10_WB.instance_to_wrap.host_row2\[85\] team_10_WB.instance_to_wrap.dispFSM.guesses\[61\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3365_ team_10_WB.instance_to_wrap.host_row2\[65\] team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload18_A clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1951__A team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3296_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ _1674_ net297 vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a31o_1
X_2316_ net225 net226 _0850_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__and3b_1
X_2247_ _0793_ net213 _0802_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] _1028_
+ vssd1 vssd1 vccd1 vccd1 _1029_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout183_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2178_ _0968_ team_10_WB.instance_to_wrap.correct\[1\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0654_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3118__A team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput46 net46 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 gpio_out[34] sky130_fd_sc_hd__buf_2
XANTENNA__4010__Q team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3358__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4322__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3150_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] _1278_ _1568_ vssd1 vssd1 vccd1
+ vccd1 _1580_ sky130_fd_sc_hd__a21o_1
X_2101_ team_10_WB.instance_to_wrap.dispFSM.guesses\[11\] net115 net136 team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__o22a_1
XANTENNA__4472__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3081_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2032_ net195 _0903_ net137 vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3050__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3983_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[20\]
+ _0051_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2934_ net602 net156 net125 net613 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[39\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2865_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\] _1454_ vssd1 vssd1
+ vccd1 vccd1 _1455_ sky130_fd_sc_hd__and2_1
X_4604_ net379 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__3349__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2541__S _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4535_ net347 vssd1 vssd1 vccd1 vccd1 DAT_O[9] sky130_fd_sc_hd__buf_2
X_2796_ _1405_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4466_ clknet_leaf_1_wb_clk_i net591 _0449_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3417_ team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] _1715_ _1791_ _1792_ vssd1
+ vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__a211o_1
X_4397_ clknet_leaf_3_wb_clk_i _0782_ _0380_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_3348_ team_10_WB.instance_to_wrap.host_row2\[64\] team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3279_ net634 _1664_ net231 vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout186_X net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3401__A net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2017__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_48_Left_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2251__B1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Left_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2214__X _1000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2650_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ _1224_ _1311_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_10_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2581_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\] _0904_ _0906_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4320_ clknet_leaf_16_wb_clk_i _0710_ _0309_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4251_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[7\]
+ _0240_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3202_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\]
+ _1392_ vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4182_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\]
+ _0171_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[44\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3133_ net220 _0905_ _1562_ _0907_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4218__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3064_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] _1526_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] sky130_fd_sc_hd__mux2_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2015_ _0887_ _0892_ net227 vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__or3b_1
XANTENNA__2536__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2490__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout146_A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[3\]
+ _0034_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4368__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2917_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\] net154 net123 net656
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[22\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3897_ net256 vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2848_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\] _1442_ vssd1 vssd1
+ vccd1 vccd1 _1444_ sky130_fd_sc_hd__and2_1
X_2779_ net728 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\] vssd1 vssd1 vccd1
+ vccd1 _1389_ sky130_fd_sc_hd__nand2_1
XANTENNA__4202__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4518_ net330 vssd1 vssd1 vccd1 vccd1 ADR_O[25] sky130_fd_sc_hd__buf_2
Xhold153 net65 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] vssd1 vssd1 vccd1
+ vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold142 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\] vssd1 vssd1 vccd1
+ vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 team_10_WB.instance_to_wrap.dispFSM.guesses\[15\] vssd1 vssd1 vccd1 vccd1
+ net577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 net70 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[6\]
+ _0432_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xhold164 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[21\] vssd1 vssd1
+ vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\] vssd1 vssd1 vccd1
+ vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1
+ vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2481__B1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4628__397 vssd1 vssd1 vccd1 vccd1 _4628__397/HI net397 sky130_fd_sc_hd__conb_1
XFILLER_0_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3016__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3820_ net254 vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3751_ net280 vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2702_ net226 net222 net300 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__mux2_1
XFILLER_0_40_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1983__C1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3682_ net248 vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2633_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] _1285_ _1290_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1300_ vssd1 vssd1 vccd1 vccd1 _0011_ sky130_fd_sc_hd__a221o_1
X_2564_ _1059_ _1250_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1
+ vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4303_ clknet_leaf_15_wb_clk_i _0693_ _0292_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2495_ net232 _1177_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_288 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4234_ clknet_leaf_21_wb_clk_i _0647_ _0223_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4040__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4165_ clknet_leaf_24_wb_clk_i _0634_ _0154_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3116_ net585 net4 _1548_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__mux2_1
X_4096_ clknet_leaf_11_wb_clk_i _0567_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3047_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__mux2_1
XANTENNA__4190__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout149_X net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3949_ clknet_leaf_23_wb_clk_i _0012_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4554__366 vssd1 vssd1 vccd1 vccd1 _4554__366/HI net366 sky130_fd_sc_hd__conb_1
XFILLER_0_56_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1980__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4063__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2280_ net219 _0952_ _1023_ _1060_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3323__X _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3803_ net272 vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] net148 vssd1 vssd1
+ vccd1 vccd1 _0884_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4497__309 vssd1 vssd1 vccd1 vccd1 _4497__309/HI net309 sky130_fd_sc_hd__conb_1
X_3734_ net293 vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3665_ net278 vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__inv_2
XANTENNA__4406__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1956__C1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2616_ _0015_ _0012_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3596_ net275 vssd1 vssd1 vccd1 vccd1 _0128_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2547_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _1239_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_54_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2478_ net528 net129 _1189_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\]
+ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__o22a_1
X_4217_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[79\]
+ _0206_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[79\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3476__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4148_ clknet_leaf_11_wb_clk_i _0619_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout266_X net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4079_ clknet_leaf_21_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[10\]
+ _0099_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2987__B2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4086__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1864__A team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 net266 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout282 net283 vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout271 net272 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__buf_4
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__buf_4
XFILLER_0_9_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4643__412 vssd1 vssd1 vccd1 vccd1 _4643__412/HI net412 sky130_fd_sc_hd__conb_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2978__B2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2206__Y _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4429__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3465__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3450_ _1781_ _1820_ _1824_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3381_ team_10_WB.instance_to_wrap.host_row1\[58\] team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1759_ sky130_fd_sc_hd__mux2_1
X_2401_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ _1160_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2332_ _0843_ net196 _0810_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2263_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0800_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ _0790_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a221o_1
X_4002_ clknet_leaf_24_wb_clk_i _0490_ net270 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3458__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2194_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] _0801_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ _0795_ _0982_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2969__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2544__S _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2969__B2 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1978_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] net150 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3717_ net236 vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3648_ net254 vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_3579_ net262 vssd1 vssd1 vccd1 vccd1 _0111_ sky130_fd_sc_hd__inv_2
XANTENNA__3946__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold13 team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] vssd1 vssd1 vccd1 vccd1 net470
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1
+ net503 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
Xhold35 team_10_WB.instance_to_wrap.message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1
+ net492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] vssd1 vssd1 vccd1 vccd1 net481
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\] vssd1 vssd1 vccd1 vccd1
+ net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] vssd1 vssd1 vccd1 vccd1
+ net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 team_10_WB.instance_to_wrap.host_row1\[47\] vssd1 vssd1 vccd1 vccd1 net525
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4008__Q team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3082__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2896__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4101__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload4_A clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3073__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2950_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\] net165 _1478_ net216 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[2\] sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_33_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _0825_ sky130_fd_sc_hd__inv_2
X_2881_ net193 _1464_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[3\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4620_ net392 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_38_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4551_ net363 vssd1 vssd1 vccd1 vccd1 DAT_O[25] sky130_fd_sc_hd__buf_2
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3969__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3502_ net250 vssd1 vssd1 vccd1 vccd1 _0034_ sky130_fd_sc_hd__inv_2
X_4482_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[39\]
+ _0465_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3433_ team_10_WB.instance_to_wrap.host_row1\[69\] net302 _1703_ vssd1 vssd1 vccd1
+ vccd1 _1808_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3364_ _1738_ _1742_ _1736_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_27_Left_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3295_ net295 _1676_ _1677_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__nor3_1
XANTENNA__2539__S _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2315_ _0868_ _1090_ net4 vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__or3b_1
X_2246_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _0804_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__a2bb2o_1
X_2177_ _0936_ _0962_ _0967_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout131_X net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3367__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4124__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput47 net47 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4274__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2869__B1 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2100_ team_10_WB.instance_to_wrap.dispFSM.guesses\[12\] net109 net136 net682 vssd1
+ vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__o22a_1
X_3080_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] _1534_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[76\] sky130_fd_sc_hd__mux2_1
X_2031_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _0886_ _0910_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3982_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[19\]
+ _0050_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_2933_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] net154 net122 net686
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[38\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2864_ _1454_ net176 _1453_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[8\]
+ sky130_fd_sc_hd__and3b_1
X_4603_ net378 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_2795_ net230 _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4534_ net346 vssd1 vssd1 vccd1 vccd1 DAT_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_29_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4465_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[22\]
+ _0448_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload30_A clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4297__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4396_ clknet_leaf_6_wb_clk_i _0781_ _0379_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\]
+ sky130_fd_sc_hd__dfstp_2
X_3416_ team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] net171 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3347_ _1682_ _1686_ _1688_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__and3_1
X_3278_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\]
+ _1663_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout179_X net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2229_ team_10_WB.instance_to_wrap.message_reg.state\[0\] net145 _0807_ vssd1 vssd1
+ vccd1 vccd1 _0647_ sky130_fd_sc_hd__o21a_1
XANTENNA__3401__B net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2017__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input21_A wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2580_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\] _0906_ _1262_ _1263_
+ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_231 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[6\]
+ _0239_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3201_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\]
+ _1391_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1
+ _1618_ sky130_fd_sc_hd__a31o_1
X_4181_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\]
+ _0170_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[43\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3132_ _0890_ _0899_ _1259_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__or3_1
X_3063_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2014_ net2 net3 net4 net5 net300 vssd1 vssd1 vccd1 vccd1 _0897_ sky130_fd_sc_hd__o41a_1
XFILLER_0_54_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3965_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[2\]
+ _0033_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3896_ net256 vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__inv_2
X_2916_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\] _1181_ _1472_ net620
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[21\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__3945__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2847_ _1442_ _1443_ net176 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\] vssd1 vssd1 vccd1
+ vccd1 net567 sky130_fd_sc_hd__dlygate4sd3_1
X_2778_ net464 _1388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[29\]
+ sky130_fd_sc_hd__xor2_1
X_4517_ net329 vssd1 vssd1 vccd1 vccd1 ADR_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold132 team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] vssd1 vssd1 vccd1 vccd1
+ net589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] vssd1 vssd1 vccd1
+ vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _0682_ vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\] vssd1 vssd1 vccd1
+ vccd1 net622 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] vssd1 vssd1 vccd1 vccd1
+ net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4448_ clknet_leaf_27_wb_clk_i net495 _0431_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold154 team_10_WB.instance_to_wrap.dispFSM.guesses\[71\] vssd1 vssd1 vccd1 vccd1
+ net611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] vssd1 vssd1 vccd1
+ vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] vssd1 vssd1 vccd1 vccd1
+ net644 sky130_fd_sc_hd__dlygate4sd3_1
X_4379_ clknet_leaf_6_wb_clk_i _0764_ _0362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_42_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2233__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4462__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3249__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_654 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3750_ net296 vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_41_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_816 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2701_ team_10_WB.instance_to_wrap.host_col\[0\] net223 net300 vssd1 vssd1 vccd1
+ vccd1 net78 sky130_fd_sc_hd__mux2_1
XFILLER_0_27_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3681_ net279 vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2632_ net195 _1281_ _1298_ _0903_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2563_ net219 _0948_ net134 vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3056__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4302_ clknet_leaf_17_wb_clk_i _0692_ _0291_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2494_ net515 net130 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] vssd1
+ vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__a22o_1
X_4233_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[2\]
+ _0222_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4164_ clknet_leaf_28_wb_clk_i _0633_ _0153_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4095_ clknet_leaf_12_wb_clk_i _0566_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3115_ net547 net3 _1548_ vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__mux2_1
X_3046_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _1517_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[59\] sky130_fd_sc_hd__mux2_1
XANTENNA__4335__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2463__B2 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2463__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4660__429 vssd1 vssd1 vccd1 vccd1 _4660__429/HI net429 sky130_fd_sc_hd__conb_1
XANTENNA__3412__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3948_ clknet_leaf_21_wb_clk_i _0011_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1974__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3879_ net275 vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4669__432 vssd1 vssd1 vccd1 vccd1 _4669__432/HI net432 sky130_fd_sc_hd__conb_1
X_4565__441 vssd1 vssd1 vccd1 vccd1 net441 _4565__441/LO sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_1_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4208__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2221__A _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4358__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3802_ net292 vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__inv_2
X_1994_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] net148 net118
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1 vccd1 _0754_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3733_ net237 vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3664_ net268 vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload30 clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__inv_6
X_2615_ _1270_ _1282_ _1293_ _1275_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0012_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2131__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ net253 vssd1 vssd1 vccd1 vccd1 _0127_ sky130_fd_sc_hd__inv_2
X_2546_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_54_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2477_ net552 net131 _1185_ _1212_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__a22o_1
X_4216_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[78\]
+ _0205_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[78\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4147_ clknet_leaf_13_wb_clk_i _0618_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__dfxtp_1
X_4588__452 vssd1 vssd1 vccd1 vccd1 net452 _4588__452/LO sky130_fd_sc_hd__conb_1
X_4078_ clknet_leaf_21_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[9\]
+ _0098_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3029_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__mux2_1
XANTENNA__2436__B2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload2 clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
X_4521__333 vssd1 vssd1 vccd1 vccd1 _4521__333/HI net333 sky130_fd_sc_hd__conb_1
XFILLER_0_34_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2911__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1880__A team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 net252 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__buf_4
Xfanout283 net299 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__buf_2
Xfanout261 net262 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_4
Xfanout272 net274 vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2124__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout294 net298 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4030__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4180__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2400_ team_10_WB.instance_to_wrap.clock_div.count\[11\] _1161_ _1162_ team_10_WB.instance_to_wrap.clock_div.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3380_ _1754_ _1755_ _1757_ vssd1 vssd1 vccd1 vccd1 _1758_ sky130_fd_sc_hd__or3_1
XFILLER_0_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2331_ _0844_ net196 _0809_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__a21o_1
XANTENNA__2902__A2 _1181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3481__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2262_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] net216 vssd1 vssd1 vccd1
+ vccd1 _1044_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4001_ clknet_leaf_24_wb_clk_i _0489_ net270 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2193_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] _0804_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__o22a_1
XANTENNA__2969__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4505__317 vssd1 vssd1 vccd1 vccd1 _4505__317/HI net317 sky130_fd_sc_hd__conb_1
XFILLER_0_8_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1977_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] net146 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[20\]
+ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout121_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3716_ net240 vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ net258 vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3578_ net263 vssd1 vssd1 vccd1 vccd1 _0110_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2529_ net465 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0512_ sky130_fd_sc_hd__mux2_1
Xhold14 _0508_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 team_10_WB.instance_to_wrap.host_row1\[42\] vssd1 vssd1 vccd1 vccd1 net504
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 team_10_WB.instance_to_wrap.host_row1\[64\] vssd1 vssd1 vccd1 vccd1 net493
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 _0507_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 team_10_WB.instance_to_wrap.host_row1\[40\] vssd1 vssd1 vccd1 vccd1 net515
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\] vssd1 vssd1 vccd1
+ vccd1 net526 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4053__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3385__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1875__A team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1900_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1 vssd1 vccd1 vccd1
+ _0824_ sky130_fd_sc_hd__inv_2
X_2880_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[3\] net1 _1463_ vssd1 vssd1 vccd1
+ vccd1 _1464_ sky130_fd_sc_hd__mux2_1
XANTENNA__3376__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4550_ net362 vssd1 vssd1 vccd1 vccd1 DAT_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_53_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4481_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[38\]
+ _0464_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3501_ net250 vssd1 vssd1 vccd1 vccd1 _0033_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3432_ team_10_WB.instance_to_wrap.host_row1\[101\] net302 _1776_ _1806_ vssd1 vssd1
+ vccd1 vccd1 _1807_ sky130_fd_sc_hd__o22a_1
X_3363_ _1739_ _1740_ _1741_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3064__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3294_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\]
+ _1672_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__and3_1
X_2314_ net225 net226 _0850_ _0818_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__o211ai_1
X_2245_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _0800_ _0802_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ _1026_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__o221a_1
X_2176_ _0959_ _0960_ _0961_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4076__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout169_A _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4679_ net183 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_X clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput48 net48 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XFILLER_0_11_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4419__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3358__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2213__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2566__B1 net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2869__A1 team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4099__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ net195 _0903_ net144 vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__a21o_1
XANTENNA__2097__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3981_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[18\]
+ _0049_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2932_ net735 net156 net125 net615 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[37\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2863_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\]
+ _1450_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__and3_1
X_4602_ net377 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
X_2794_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[5\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_903 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4621__393 vssd1 vssd1 vccd1 vccd1 _4621__393/HI net393 sky130_fd_sc_hd__conb_1
X_4533_ net345 vssd1 vssd1 vccd1 vccd1 DAT_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_13_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4464_ clknet_leaf_27_wb_clk_i net621 _0447_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1962__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4395_ clknet_leaf_6_wb_clk_i _0780_ _0378_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload23_A clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3415_ team_10_WB.instance_to_wrap.dispFSM.guesses\[60\] _1701_ net168 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\]
+ _1771_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__a221o_1
X_3346_ _1722_ _1725_ _1713_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__o21a_1
X_3277_ net548 _1661_ _1665_ vssd1 vssd1 vccd1 vccd1 _0564_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2228_ net492 _1011_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_37_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2159_ _0924_ _0945_ _0951_ _0953_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__or4_1
XANTENNA__3401__C net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2984__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4391__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3959__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4212__Q team_10_WB.instance_to_wrap.host_row2\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3200_ net172 _1617_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__nor2_1
X_4180_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[42\]
+ _0169_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[42\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2894__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3131_ net221 _1259_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3062_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] _1525_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[67\] sky130_fd_sc_hd__mux2_1
XFILLER_0_54_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2013_ net301 net5 vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2490__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4114__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3964_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[1\]
+ _0032_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3895_ net277 vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__inv_2
X_2915_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\] net152 net121 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[20\]
+ sky130_fd_sc_hd__o22a_1
X_2846_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold100 team_10_WB.instance_to_wrap.host_row1\[77\] vssd1 vssd1 vccd1 vccd1 net557
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ _1387_ _1388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[28\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4516_ net328 vssd1 vssd1 vccd1 vccd1 ADR_O[23] sky130_fd_sc_hd__buf_2
Xhold144 team_10_WB.instance_to_wrap.host_row1\[65\] vssd1 vssd1 vccd1 vccd1 net601
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 team_10_WB.instance_to_wrap.host_row1\[57\] vssd1 vssd1 vccd1 vccd1 net568
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold133 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\] vssd1 vssd1 vccd1
+ vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] vssd1 vssd1 vccd1 vccd1
+ net579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\] vssd1 vssd1 vccd1 vccd1
+ net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\] vssd1 vssd1 vccd1
+ vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[4\]
+ _0430_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2950__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 team_10_WB.instance_to_wrap.clock_div.count\[28\] vssd1 vssd1 vccd1 vccd1
+ net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\] vssd1 vssd1 vccd1
+ vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold188 team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] vssd1 vssd1 vccd1 vccd1
+ net645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input6_A gpio_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4378_ clknet_leaf_1_wb_clk_i _0763_ _0361_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3329_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _1682_ _1688_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__and4_1
XANTENNA__2466__C1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2233__A2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2941__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4137__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2219__A net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1085 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3421__A1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4287__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3421__B2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_828 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2700_ _1342_ _1344_ _1238_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.tx_serial
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ net268 vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__inv_2
X_2631_ _0911_ _1298_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__nor2_1
X_2562_ net134 _0972_ _1249_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__and3_1
X_4301_ clknet_leaf_14_wb_clk_i _0691_ _0290_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[24\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2932__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2493_ net553 net133 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] vssd1
+ vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4232_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[1\]
+ _0221_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4163_ clknet_leaf_24_wb_clk_i _0632_ _0152_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4094_ clknet_leaf_12_wb_clk_i _0565_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_3114_ net520 net2 _1548_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__mux2_1
X_3045_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2463__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout151_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2416__X _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3947_ clknet_leaf_3_wb_clk_i _0479_ _0021_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1974__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3878_ net275 vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2829_ _1411_ _1418_ _1426_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__and3_1
XANTENNA__1974__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2923__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_X net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2439__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1878__A net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1094 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2914__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3801_ net292 vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] _0874_ _0883_ net158 vssd1
+ vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1956__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3732_ net238 vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__inv_2
X_3663_ net278 vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload20 clknet_leaf_23_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_15_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2614_ _0824_ _1287_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2905__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3594_ net268 vssd1 vssd1 vccd1 vccd1 _0126_ sky130_fd_sc_hd__inv_2
XANTENNA__4302__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2545_ net228 net458 _1216_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__mux2_1
XANTENNA__2381__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4400__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2476_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] net186 vssd1 vssd1 vccd1
+ vccd1 _1212_ sky130_fd_sc_hd__or2_1
X_4215_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[77\]
+ _0204_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[77\] sky130_fd_sc_hd__dfrtp_1
X_4146_ clknet_leaf_11_wb_clk_i _0617_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.lcd_rs
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout199_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4452__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4077_ clknet_leaf_21_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[8\]
+ _0097_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3028_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] _1508_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[50\] sky130_fd_sc_hd__mux2_1
XFILLER_0_47_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_143 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4560__372 vssd1 vssd1 vccd1 vccd1 _4560__372/HI net372 sky130_fd_sc_hd__conb_1
Xclkload3 clknet_leaf_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload3/Y sky130_fd_sc_hd__inv_8
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout240 net241 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_4
Xfanout262 net265 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 net252 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_4
Xfanout273 net274 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
Xfanout295 net297 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_4
Xfanout284 net288 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_17_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3388__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4325__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4220__Q team_10_WB.instance_to_wrap.host_row2\[82\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2330_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] _0819_ _0849_ vssd1
+ vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__or3_1
XANTENNA__4475__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2261_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] _0799_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ _1042_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__a221o_1
XANTENNA__3312__B1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ clknet_leaf_24_wb_clk_i _0488_ net270 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2192_ team_10_WB.instance_to_wrap.gamelogic.setWord\[11\] _0802_ _0804_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_47_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4544__356 vssd1 vssd1 vccd1 vccd1 _4544__356/HI net356 sky130_fd_sc_hd__conb_1
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3379__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1976_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] _0874_ _0880_ net159 vssd1
+ vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3715_ net240 vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1965__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout114_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ net256 vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
XANTENNA__4017__RESET_B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ net271 vssd1 vssd1 vccd1 vccd1 _0109_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2528_ _1233_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold15 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] vssd1 vssd1 vccd1 vccd1 net472
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\] vssd1 vssd1 vccd1 vccd1
+ net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 team_10_WB.instance_to_wrap.message_reg.msg\[5\] vssd1 vssd1 vccd1 vccd1 net483
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] net197 _1185_
+ _1202_ net132 vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a221o_1
Xhold48 team_10_WB.instance_to_wrap.host_row1\[71\] vssd1 vssd1 vccd1 vccd1 net505
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold59 team_10_WB.instance_to_wrap.host_row1\[63\] vssd1 vssd1 vccd1 vccd1 net516
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4129_ clknet_leaf_18_wb_clk_i _0600_ _0128_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[64\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3992__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4348__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3500_ net251 vssd1 vssd1 vccd1 vccd1 _0032_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4480_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[37\]
+ _0463_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_3431_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1805_ _1686_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3362_ team_10_WB.instance_to_wrap.host_row2\[49\] net170 _1708_ team_10_WB.instance_to_wrap.host_row1\[73\]
+ vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ net229 _0848_ net196 net225 vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3293_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\] _1674_ vssd1 vssd1 vccd1
+ vccd1 _1676_ sky130_fd_sc_hd__nor2_1
X_2244_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0798_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_10_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2175_ _0966_ team_10_WB.instance_to_wrap.correct\[2\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0655_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2137__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1959_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] net146 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[34\]
+ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4678_ net434 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[17] sky130_fd_sc_hd__buf_2
XANTENNA_fanout117_X net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3629_ net253 vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__inv_2
X_4633__402 vssd1 vssd1 vccd1 vccd1 _4633__402/HI net402 sky130_fd_sc_hd__conb_1
Xoutput49 net49 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_8_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4170__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2263__B1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3460__C1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2869__A2 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[17\]
+ _0048_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2931_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] net151 net121 net653
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[36\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3451__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4601_ net376 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2862_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ _1448_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[8\] vssd1 vssd1 vccd1
+ vccd1 _1453_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2793_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] _1393_ _1395_ _1402_
+ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__or4_4
XFILLER_0_41_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4532_ net344 vssd1 vssd1 vccd1 vccd1 DAT_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4463_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[20\]
+ _0446_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3414_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1704_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[68\]
+ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2420__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4394_ clknet_leaf_1_wb_clk_i _0779_ _0377_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[31\]
+ sky130_fd_sc_hd__dfrtp_2
X_3345_ _1716_ _1723_ _1724_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__or3_1
XANTENNA_clkload16_A clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3276_ net295 _1664_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nor2_1
X_2227_ team_10_WB.instance_to_wrap.uart_transmitter.state\[1\] _1009_ _1010_ _0808_
+ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__o22a_1
XANTENNA__2419__X _1181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4193__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2493__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2158_ net219 net218 _0947_ _0952_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2089_ net573 net145 net108 net592 vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2984__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2236__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_3__f_wb_clk_i_X clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3130_ _1286_ _1554_ _1560_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3061_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Left_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2475__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2012_ net301 net5 vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[0\]
+ _0031_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_3894_ net260 vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__inv_2
X_2914_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\] net153 net121 net719
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[19\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4409__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2845_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1442_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1986__C1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4515_ net327 vssd1 vssd1 vccd1 vccd1 ADR_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_5_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2776_ team_10_WB.instance_to_wrap.clock_div.count\[27\] team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ team_10_WB.instance_to_wrap.clock_div.count\[28\] _1384_ vssd1 vssd1 vccd1 vccd1
+ _1388_ sky130_fd_sc_hd__and4_1
Xhold101 team_10_WB.instance_to_wrap.dispFSM.guesses\[47\] vssd1 vssd1 vccd1 vccd1
+ net558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 team_10_WB.instance_to_wrap.clock_div.count\[1\] vssd1 vssd1 vccd1 vccd1
+ net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[23\] vssd1 vssd1
+ vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 team_10_WB.instance_to_wrap.dispFSM.guesses\[61\] vssd1 vssd1 vccd1 vccd1
+ net569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\] vssd1 vssd1 vccd1 vccd1
+ net624 sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[3\]
+ _0429_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2950__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2150__A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold145 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[47\] vssd1 vssd1 vccd1
+ vccd1 net602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[39\] vssd1 vssd1 vccd1
+ vccd1 net613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\] vssd1 vssd1 vccd1 vccd1
+ net635 sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ clknet_leaf_7_wb_clk_i _0762_ _0360_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\]
+ sky130_fd_sc_hd__dfstp_2
Xhold189 team_10_WB.instance_to_wrap.dispFSM.guesses\[43\] vssd1 vssd1 vccd1 vccd1
+ net646 sky130_fd_sc_hd__dlygate4sd3_1
X_3328_ _1697_ _1707_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__nor2_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3259_ net296 _1653_ vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout184_X net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2466__B1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2941__A1 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1097 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2630_ _0886_ _0909_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__nor2_1
XANTENNA__1983__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3337__Y _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2561_ net219 net218 _0947_ _1034_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__a41o_1
X_2492_ net504 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\] vssd1
+ vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__a22o_1
X_4300_ clknet_leaf_19_wb_clk_i _0690_ _0289_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4231_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_state\[0\]
+ _0220_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_4162_ clknet_leaf_24_wb_clk_i _0631_ _0151_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4093_ clknet_leaf_12_wb_clk_i _0564_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3113_ net560 net220 _1548_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__mux2_1
XANTENNA__2448__B1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3044_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] _1516_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[58\] sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_X clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2999__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout144_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ clknet_leaf_1_wb_clk_i _0478_ _0020_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__3412__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1974__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3877_ net253 vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__inv_2
X_2828_ _1409_ _0513_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__nand2_1
XANTENNA__4381__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2759_ team_10_WB.instance_to_wrap.clock_div.count\[21\] _1376_ vssd1 vssd1 vccd1
+ vccd1 _1378_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4429_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[26\]
+ _0412_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3479__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2439__B1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3167__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4104__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3800_ net293 vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3731_ net237 vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__inv_2
X_1992_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] net149 vssd1 vssd1
+ vccd1 vccd1 _0883_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3662_ net257 vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__inv_2
Xclkload10 clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload10/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1956__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2613_ _0016_ _0014_ _0015_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
Xclkload21 clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__inv_6
X_3593_ net253 vssd1 vssd1 vccd1 vccd1 _0125_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2544_ team_10_WB.instance_to_wrap.host_col\[0\] _1237_ _1179_ vssd1 vssd1 vccd1
+ vccd1 _0484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2475_ net507 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\]
+ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__a22o_1
X_4214_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[76\]
+ _0203_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[76\] sky130_fd_sc_hd__dfrtp_1
X_4145_ clknet_leaf_17_wb_clk_i _0616_ _0144_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[101\]
+ sky130_fd_sc_hd__dfrtp_1
X_4076_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[7\]
+ _0096_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3027_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout147_X net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3929_ net240 vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload4 clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1920__A_N net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4127__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _0018_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xfanout241 net243 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__buf_4
XANTENNA__4277__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net265 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_4
Xfanout274 net283 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 net255 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_2
Xfanout296 net297 vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_4
Xfanout285 net287 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2232__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2899__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4650__419 vssd1 vssd1 vccd1 vccd1 _4650__419/HI net419 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_53_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2260_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0800_ vssd1 vssd1 vccd1
+ vccd1 _1042_ sky130_fd_sc_hd__nor2_1
X_2191_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] team_10_WB.instance_to_wrap.gamelogic.letter\[5\]
+ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1975_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] net148 vssd1 vssd1 vccd1
+ vccd1 _0880_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3714_ net236 vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3645_ net256 vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3576_ net264 vssd1 vssd1 vccd1 vccd1 _0108_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2527_ team_10_WB.instance_to_wrap.uart_receiver.state\[0\] team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] vssd1 vssd1 vccd1 vccd1 _1233_
+ sky130_fd_sc_hd__or3b_4
X_2458_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] net186 vssd1 vssd1 vccd1
+ vccd1 _1202_ sky130_fd_sc_hd__or2_1
Xhold38 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[5\] vssd1 vssd1 vccd1
+ vccd1 net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 _0509_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 team_10_WB.instance_to_wrap.dispFSM.guesses\[5\] vssd1 vssd1 vccd1 vccd1 net484
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_3_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2389_ _0844_ net587 _1158_ vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__mux2_1
Xhold49 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[10\] vssd1 vssd1 vccd1
+ vccd1 net506 sky130_fd_sc_hd__dlygate4sd3_1
X_4128_ clknet_leaf_26_wb_clk_i _0599_ _0127_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3067__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4059_ clknet_leaf_15_wb_clk_i _0544_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input37_A wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3058__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3103__S net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4442__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ net210 _0817_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3361_ team_10_WB.instance_to_wrap.host_row1\[49\] _1699_ net169 team_10_WB.instance_to_wrap.host_row1\[57\]
+ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2312_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__inv_2
X_3292_ net536 _1672_ _1675_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2243_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] _0805_ vssd1 vssd1 vccd1
+ vccd1 _1025_ sky130_fd_sc_hd__or2_1
X_4511__323 vssd1 vssd1 vccd1 vccd1 _4511__323/HI net323 sky130_fd_sc_hd__conb_1
X_2174_ _0964_ _0965_ vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2424__Y _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1958_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[35\]
+ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4677_ net183 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_1
X_1889_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\] vssd1 vssd1 vccd1 vccd1
+ _0813_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3628_ net268 vssd1 vssd1 vccd1 vccd1 _0160_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3559_ net289 vssd1 vssd1 vccd1 vccd1 _0091_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3288__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3712__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2263__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3460__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4465__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2998__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2213__D net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3279__B1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3622__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload2_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4226__Q team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2930_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] net151 net120 net673
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[35\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4600_ net457 vssd1 vssd1 vccd1 vccd1 gpio_oeb[37] sky130_fd_sc_hd__buf_2
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ net527 _1450_ _1452_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_2792_ _1396_ _1400_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4531_ net343 vssd1 vssd1 vccd1 vccd1 DAT_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4656__425 vssd1 vssd1 vccd1 vccd1 _4656__425/HI net425 sky130_fd_sc_hd__conb_1
X_4462_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[19\]
+ _0445_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_13_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3413_ team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] net181 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4393_ clknet_leaf_7_wb_clk_i _0778_ _0376_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2420__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3344_ team_10_WB.instance_to_wrap.dispFSM.guesses\[0\] _1717_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[64\]
+ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__a22o_1
X_3275_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] _1661_ vssd1 vssd1 vccd1
+ vccd1 _1664_ sky130_fd_sc_hd__and2_1
X_2226_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] vssd1 vssd1 vccd1 vccd1
+ _1010_ sky130_fd_sc_hd__or3b_1
XANTENNA__4338__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ net218 _0916_ vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2088_ team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] net114 net141 net733 vssd1
+ vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4488__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4600__457 vssd1 vssd1 vccd1 vccd1 net457 _4600__457/LO sky130_fd_sc_hd__conb_1
XFILLER_0_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3433__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3617__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output68_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] _1524_ net203 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[66\] sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_12_wb_clk_i_X clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2011_ net301 net4 vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3424__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ clknet_leaf_21_wb_clk_i _0482_ _0030_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3893_ net262 vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__inv_2
X_2913_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\] net151 net120 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[18\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2844_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net490 _1441_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4010__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514_ net326 vssd1 vssd1 vccd1 vccd1 ADR_O[21] sky130_fd_sc_hd__buf_2
XANTENNA__2431__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2775_ team_10_WB.instance_to_wrap.clock_div.count\[27\] _1386_ net623 vssd1 vssd1
+ vccd1 vccd1 _1387_ sky130_fd_sc_hd__a21oi_1
Xhold124 team_10_WB.instance_to_wrap.host_row1\[70\] vssd1 vssd1 vccd1 vccd1 net581
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] vssd1 vssd1 vccd1 vccd1
+ net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _0728_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _0714_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4445_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[2\]
+ _0428_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
Xhold146 team_10_WB.instance_to_wrap.clock_div.count\[24\] vssd1 vssd1 vccd1 vccd1
+ net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\] vssd1 vssd1 vccd1
+ vccd1 net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 team_10_WB.instance_to_wrap.host_row1\[60\] vssd1 vssd1 vccd1 vccd1 net614
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\] vssd1 vssd1 vccd1 vccd1
+ net636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4160__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4376_ clknet_leaf_27_wb_clk_i _0761_ _0359_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__3360__C1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3327_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _1707_ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout291_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3258_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] _1651_ vssd1 vssd1 vccd1
+ vccd1 _1653_ sky130_fd_sc_hd__and2_1
X_3189_ net298 net178 _1610_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout177_X net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2466__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2209_ net487 _0996_ _0992_ vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3415__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1977__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3351__C1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4033__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4183__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2560_ _0973_ _1248_ vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2491_ net538 net133 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] vssd1
+ vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__a22o_1
XANTENNA__2932__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4230_ clknet_leaf_0_wb_clk_i _0646_ _0219_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4161_ clknet_leaf_28_wb_clk_i _0630_ _0150_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4092_ clknet_leaf_13_wb_clk_i _0563_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_3112_ net542 net221 _1548_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__mux2_1
X_3043_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2426__A _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3945_ clknet_leaf_3_wb_clk_i _0477_ _0019_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1959__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3876_ net267 vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2827_ _1407_ _1418_ _1429_ _1427_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2758_ team_10_WB.instance_to_wrap.clock_div.count\[21\] _1376_ vssd1 vssd1 vccd1
+ vccd1 _1377_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout304_A net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4428_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[25\]
+ _0411_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2689_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] _1336_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_18_Left_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2136__A0 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4359_ clknet_leaf_10_wb_clk_i _0002_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4056__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3720__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Left_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2914__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Left_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4572__448 vssd1 vssd1 vccd1 vccd1 net448 _4572__448/LO sky130_fd_sc_hd__conb_1
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1991_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] net149 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3730_ net236 vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3661_ net256 vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__inv_2
Xclkload11 clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__inv_8
X_2612_ net195 _0909_ _1292_ _1290_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0015_ sky130_fd_sc_hd__a32o_1
Xclkload22 clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_24_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3592_ net268 vssd1 vssd1 vccd1 vccd1 _0124_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2905__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2543_ _0819_ team_10_WB.instance_to_wrap.host_col\[0\] _0851_ vssd1 vssd1 vccd1
+ vccd1 _1237_ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2474_ net523 net129 _1211_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__o21a_1
X_4213_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[75\]
+ _0202_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[75\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__4079__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4144_ clknet_leaf_2_wb_clk_i _0615_ _0143_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_4075_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[6\]
+ _0095_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3026_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _1507_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[49\] sky130_fd_sc_hd__mux2_1
XANTENNA__3094__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3397__A2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ net240 vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__inv_2
Xclkload5 clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload5/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_61_435 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3859_ net261 vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout231 _0018_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_2
Xfanout220 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] vssd1 vssd1 vccd1
+ vccd1 net220 sky130_fd_sc_hd__buf_2
Xfanout242 net243 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_4
Xfanout264 net265 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_4
Xfanout253 net255 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout297 net298 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__clkbuf_2
Xfanout275 net279 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__buf_4
Xfanout286 net287 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3388__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2190_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net213 vssd1 vssd1 vccd1
+ vccd1 _0979_ sky130_fd_sc_hd__or2_1
XANTENNA__4371__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1974_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\]
+ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__o22a_1
XANTENNA__3379__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2423__B net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3713_ net233 vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__inv_2
X_3644_ net277 vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3000__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3575_ net276 vssd1 vssd1 vccd1 vccd1 _0107_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3535__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2526_ net488 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1
+ vccd1 vccd1 _0519_ sky130_fd_sc_hd__a22o_1
X_2457_ net516 net129 _1201_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold28 _0672_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 team_10_WB.instance_to_wrap.host_row1\[61\] vssd1 vssd1 vccd1 vccd1 net474
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2388_ net5 net606 _1158_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__mux2_1
Xhold39 team_10_WB.instance_to_wrap.message_reg.msg\[4\] vssd1 vssd1 vccd1 vccd1 net496
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4127_ clknet_leaf_26_wb_clk_i _0598_ _0126_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[62\]
+ sky130_fd_sc_hd__dfrtp_1
X_4058_ clknet_leaf_15_wb_clk_i _0543_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_3009_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] net191 vssd1 vssd1 vccd1
+ vccd1 _1499_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4394__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_733 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3360_ team_10_WB.instance_to_wrap.host_row2\[57\] net180 net167 team_10_WB.instance_to_wrap.host_row2\[73\]
+ net304 vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2311_ _0841_ _1069_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__or3b_2
X_3291_ net282 _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2242_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__inv_2
X_4550__362 vssd1 vssd1 vccd1 vccd1 _4550__362/HI net362 sky130_fd_sc_hd__conb_1
X_2173_ _0959_ _0962_ _0963_ _0937_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a31o_1
XANTENNA__4117__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2418__B _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2272__A2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1957_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4676_ net183 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1888_ net220 vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout217_A team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1992__B net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_874 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3627_ net268 vssd1 vssd1 vccd1 vccd1 _0159_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3558_ net289 vssd1 vssd1 vccd1 vccd1 _0090_ sky130_fd_sc_hd__inv_2
XANTENNA__2416__A_N _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2509_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] net224 _1225_ vssd1
+ vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__and3_1
X_3489_ net241 vssd1 vssd1 vccd1 vccd1 _0021_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2263__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4493__305 vssd1 vssd1 vccd1 vccd1 _4493__305/HI net305 sky130_fd_sc_hd__conb_1
XANTENNA__3903__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4534__346 vssd1 vssd1 vccd1 vccd1 _4534__346/HI net346 sky130_fd_sc_hd__conb_1
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2860_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] _1450_ net176
+ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_26_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2791_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4530_ net342 vssd1 vssd1 vccd1 vccd1 DAT_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_13_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4461_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[18\]
+ _0444_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3412_ team_10_WB.instance_to_wrap.host_row1\[60\] net169 _1708_ team_10_WB.instance_to_wrap.host_row1\[76\]
+ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4392_ clknet_leaf_27_wb_clk_i _0777_ _0375_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_3343_ team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] net170 _1704_ team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ net232 vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__a221o_1
X_3274_ net498 _1660_ _1662_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__o21a_1
X_2225_ _0808_ team_10_WB.instance_to_wrap.uart_transmitter.state\[2\] team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__or3b_1
XANTENNA__3024__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _0949_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2087_ team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] net109 net135 net705 vssd1
+ vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2245__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\] net161 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[27\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout122_X net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_202 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4659_ net428 vssd1 vssd1 vccd1 vccd1 la_data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3723__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4432__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2236__A2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_32_Left_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2010_ net220 net221 net222 net223 vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__or4_1
XANTENNA__2475__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_46_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_X clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ clknet_leaf_21_wb_clk_i _0481_ _0029_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_63_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2912_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\] net154 net123 net676
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[17\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_63_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3892_ net265 vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2843_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ net176 vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o21ai_1
X_2774_ net532 _1386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[27\]
+ sky130_fd_sc_hd__xor2_1
X_4513_ net325 vssd1 vssd1 vccd1 vccd1 ADR_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__2935__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4305__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 team_10_WB.instance_to_wrap.clock_div.count\[13\] vssd1 vssd1 vccd1 vccd1
+ net571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\] vssd1 vssd1 vccd1 vccd1
+ net582 sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[1\]
+ _0427_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
Xhold147 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\] vssd1 vssd1 vccd1
+ vccd1 net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 team_10_WB.instance_to_wrap.host_row1\[66\] vssd1 vssd1 vccd1 vccd1 net593
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[37\] vssd1 vssd1 vccd1
+ vccd1 net615 sky130_fd_sc_hd__dlygate4sd3_1
X_4375_ clknet_leaf_8_wb_clk_i _0760_ _0358_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkload21_A clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold169 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1 vccd1
+ vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3360__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3326_ team_10_WB.instance_to_wrap.host_row2\[80\] net173 net170 team_10_WB.instance_to_wrap.host_row2\[48\]
+ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3543__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4455__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3257_ _1651_ _1652_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout284_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3188_ net298 net178 _1610_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nor3_2
XANTENNA__2466__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2208_ _0946_ _0995_ _0990_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__o21a_1
X_2139_ net134 _0934_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3718__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2926__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_728 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3103__A0 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2457__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input12_A wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3406__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3972__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4499__311 vssd1 vssd1 vccd1 vccd1 _4499__311/HI net311 sky130_fd_sc_hd__conb_1
XFILLER_0_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2490_ net529 net130 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] vssd1
+ vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_739 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3342__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4160_ clknet_leaf_24_wb_clk_i _0629_ _0149_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3111_ net522 net222 _1548_ vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__mux2_1
X_4091_ clknet_leaf_13_wb_clk_i _0562_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_3042_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] _1515_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[57\] sky130_fd_sc_hd__mux2_1
XANTENNA__2448__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ clknet_leaf_3_wb_clk_i _0476_ _0018_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3875_ net255 vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2826_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__inv_2
XANTENNA__3538__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2757_ _1375_ _1376_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[20\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2688_ _1336_ _1337_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[9\]
+ sky130_fd_sc_hd__nor2_1
X_4427_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[24\]
+ _0410_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\]
+ sky130_fd_sc_hd__dfstp_1
X_4358_ clknet_leaf_11_wb_clk_i _0001_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_input4_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4289_ clknet_leaf_12_wb_clk_i _0679_ _0278_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_3309_ _0815_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1679_ vssd1 vssd1
+ vccd1 vccd1 _1690_ sky130_fd_sc_hd__and3_1
XANTENNA__2439__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3995__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_146 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2375__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3911__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4000__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4150__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1990_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ net278 vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload23 clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__bufinv_16
Xclkload12 clknet_leaf_4_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__inv_12
X_3591_ net276 vssd1 vssd1 vccd1 vccd1 _0123_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2611_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ _1291_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_58_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2542_ net226 _1068_ _1179_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__mux2_1
XANTENNA__2366__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4212_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[74\]
+ _0201_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[74\] sky130_fd_sc_hd__dfrtp_1
X_2473_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] net198 _1185_
+ _1210_ net132 vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__a221o_1
X_4143_ clknet_leaf_8_wb_clk_i _0614_ _0142_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_4074_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[5\]
+ _0094_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3025_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout247_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ net263 vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__inv_2
X_3858_ net258 vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload6 clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__inv_4
XFILLER_0_11_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2809_ net230 _1414_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3789_ net272 vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout202_X net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout210 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1
+ vccd1 net210 sky130_fd_sc_hd__buf_2
Xfanout232 _0821_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__buf_4
Xfanout221 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] vssd1 vssd1 vccd1
+ vccd1 net221 sky130_fd_sc_hd__buf_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__buf_2
XANTENNA_input7_X net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 net255 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
Xfanout298 net299 vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_4
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4173__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2045__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2899__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2520__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2257__A team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1973_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0874_ _0879_ net157 vssd1
+ vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4624__394 vssd1 vssd1 vccd1 vccd1 _4624__394/HI net394 sky130_fd_sc_hd__conb_1
XFILLER_0_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3712_ net298 vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3643_ net264 vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4046__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3574_ net262 vssd1 vssd1 vccd1 vccd1 _0106_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3027__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2525_ net521 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1
+ vccd1 vccd1 _0520_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_5 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2456_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] net197 team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\]
+ net127 net131 vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__a221o_1
Xhold18 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] vssd1 vssd1 vccd1 vccd1
+ net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 team_10_WB.instance_to_wrap.host_row1\[62\] vssd1 vssd1 vccd1 vccd1 net486
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4196__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2387_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0856_ vssd1 vssd1 vccd1
+ vccd1 _1158_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_3_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4126_ clknet_leaf_26_wb_clk_i _0597_ _0125_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4057_ clknet_leaf_15_wb_clk_i _0542_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_3008_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\] net185 _1498_ net206
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[40\] sky130_fd_sc_hd__o211a_1
XANTENNA__3472__C1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4069__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3290_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] _1668_ vssd1 vssd1 vccd1 vccd1
+ _1674_ sky130_fd_sc_hd__and4_1
X_2310_ team_10_WB.instance_to_wrap.host_col\[0\] _0859_ _0864_ vssd1 vssd1 vccd1
+ vccd1 _1086_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2241_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] _1022_ _1013_ _1015_
+ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__or4b_2
X_2172_ _0959_ _0962_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1956_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] _0874_ _0876_ net157 vssd1
+ vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4675_ net433 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[14] sky130_fd_sc_hd__buf_2
X_1887_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 _0811_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_886 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3626_ net268 vssd1 vssd1 vccd1 vccd1 _0158_ sky130_fd_sc_hd__inv_2
XANTENNA__2980__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout112_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3557_ net289 vssd1 vssd1 vccd1 vccd1 _0089_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2508_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] _1224_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__o21a_2
X_3488_ net237 vssd1 vssd1 vccd1 vccd1 _0020_ sky130_fd_sc_hd__inv_2
X_2439_ team_10_WB.instance_to_wrap.host_row1\[74\] net132 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__a221o_1
X_4109_ clknet_leaf_8_wb_clk_i _0580_ _0108_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3460__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640__409 vssd1 vssd1 vccd1 vccd1 _4640__409/HI net409 sky130_fd_sc_hd__conb_1
XANTENNA__4211__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4361__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A wbs_stb_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2487__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3436__C1 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2254__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4460_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[17\]
+ _0443_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2270__A team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2962__B2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4391_ clknet_leaf_6_wb_clk_i _0776_ _0374_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ sky130_fd_sc_hd__dfstp_1
X_3411_ team_10_WB.instance_to_wrap.host_row2\[52\] net170 _1784_ _1786_ vssd1 vssd1
+ vccd1 vccd1 _1787_ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3342_ team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] net174 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3273_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ vssd1 vssd1 vccd1 vccd1
+ _1663_ sky130_fd_sc_hd__and4_1
X_2224_ net649 net41 _1008_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__mux2_1
XANTENNA__2478__B1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2155_ _0935_ _0948_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2086_ team_10_WB.instance_to_wrap.dispFSM.guesses\[26\] net114 net142 net650 vssd1
+ vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o22a_1
XANTENNA__4234__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4384__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2988_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\] net160 _1491_ net216
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1939_ team_10_WB.instance_to_wrap.host_message_reg.Cstate team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] _0861_ vssd1 vssd1 vccd1 vccd1
+ _0862_ sky130_fd_sc_hd__or4_1
X_4658_ net427 vssd1 vssd1 vccd1 vccd1 la_data_out[28] sky130_fd_sc_hd__buf_2
XANTENNA_fanout115_X net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2953__A1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3609_ net276 vssd1 vssd1 vccd1 vccd1 _0141_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4589_ net453 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
X_4557__369 vssd1 vssd1 vccd1 vccd1 _4557__369/HI net369 sky130_fd_sc_hd__conb_1
XFILLER_0_3_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2469__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3433__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4501__313 vssd1 vssd1 vccd1 vccd1 _4501__313/HI net313 sky130_fd_sc_hd__conb_1
XFILLER_0_2_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4107__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3960_ clknet_leaf_21_wb_clk_i _0480_ _0028_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_2911_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\] net153 net121 net687
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[16\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3424__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3891_ net261 vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__inv_2
XANTENNA__1986__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2842_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\] net176 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_60_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2773_ _1385_ _1386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[26\]
+ sky130_fd_sc_hd__nor2_1
X_4512_ net324 vssd1 vssd1 vccd1 vccd1 ADR_O[19] sky130_fd_sc_hd__buf_2
XANTENNA__2935__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold104 team_10_WB.instance_to_wrap.host_row1\[78\] vssd1 vssd1 vccd1 vccd1 net561
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 team_10_WB.instance_to_wrap.host_row1\[67\] vssd1 vssd1 vccd1 vccd1 net572
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold126 _0736_ vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[0\]
+ _0426_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xhold148 team_10_WB.instance_to_wrap.dispFSM.guesses\[67\] vssd1 vssd1 vccd1 vccd1
+ net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\] vssd1 vssd1 vccd1
+ vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\] vssd1 vssd1 vccd1 vccd1
+ net594 sky130_fd_sc_hd__dlygate4sd3_1
X_4374_ clknet_leaf_8_wb_clk_i _0759_ _0357_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload14_A clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3325_ team_10_WB.instance_to_wrap.host_row1\[64\] _1703_ net169 team_10_WB.instance_to_wrap.host_row1\[56\]
+ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3035__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3256_ _0813_ _1650_ net296 vssd1 vssd1 vccd1 vccd1 _1652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2207_ net194 _0993_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__or2_2
X_3187_ _0814_ _1607_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__or3b_4
XANTENNA_fanout277_A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2871__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2138_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ _0926_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__mux2_1
X_2069_ team_10_WB.instance_to_wrap.dispFSM.guesses\[43\] net112 net138 net685 vssd1
+ vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3415__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3103__A1 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4646__415 vssd1 vssd1 vccd1 vccd1 _4646__415/HI net415 sky130_fd_sc_hd__conb_1
XFILLER_0_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3110_ net554 net223 _1548_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ clknet_leaf_13_wb_clk_i _0561_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3041_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3943_ net299 vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ net269 vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
X_2825_ net230 _1412_ _1417_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2756_ team_10_WB.instance_to_wrap.clock_div.count\[19\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ _1372_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2687_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] _1334_ _1319_ vssd1
+ vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__o21ai_1
XANTENNA__3554__A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4422__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4426_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[23\]
+ _0409_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2315__C_N net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4357_ clknet_leaf_10_wb_clk_i _0000_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3308_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net210 _1686_ _1688_
+ _1685_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__a41o_1
X_4288_ clknet_leaf_17_wb_clk_i _0678_ _0277_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout182_X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3239_ _1642_ _1611_ _1641_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_1_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3639__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4445__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2262__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload24 clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinv_4
Xclkload13 clknet_leaf_5_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload13/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2610_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__or2_1
X_3590_ net268 vssd1 vssd1 vccd1 vccd1 _0122_ sky130_fd_sc_hd__inv_2
X_2541_ net225 _1236_ _1179_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2472_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] net186 vssd1 vssd1 vccd1
+ vccd1 _1210_ sky130_fd_sc_hd__or2_1
X_4211_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[73\]
+ _0200_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[73\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3093__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4142_ clknet_leaf_17_wb_clk_i _0613_ _0141_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_4073_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[4\]
+ _0093_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3024_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] _1506_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[48\] sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3094__A3 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3926_ net243 vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3857_ net279 vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload7 clknet_leaf_29_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload7/Y sky130_fd_sc_hd__clkinv_8
X_2808_ net210 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[2\] _1403_ vssd1
+ vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ net286 vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2739_ _1363_ _1364_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[14\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2109__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout211 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[2\] vssd1 vssd1 vccd1
+ vccd1 net211 sky130_fd_sc_hd__dlymetal6s2s_1
X_4409_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[6\]
+ _0392_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout200 net201 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout222 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\] vssd1 vssd1 vccd1
+ vccd1 net222 sky130_fd_sc_hd__buf_2
XANTENNA__3962__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout233 net239 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_4
Xfanout244 net266 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_4
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout255 net266 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_2
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__buf_4
Xfanout299 net7 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_4
Xfanout266 net7 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
Xfanout288 net291 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4318__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4468__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3242__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_X clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2257__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2446__A1_N _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2036__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1972_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] net147 vssd1 vssd1 vccd1
+ vccd1 _0879_ sky130_fd_sc_hd__or2_1
X_4691_ net184 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_1
X_3711_ net235 vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3642_ net254 vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3573_ net278 vssd1 vssd1 vccd1 vccd1 _0105_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2524_ net497 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1
+ vccd1 vccd1 _0521_ sky130_fd_sc_hd__a22o_1
X_2455_ net493 net132 _1185_ _1200_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a22o_1
X_2386_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] _1084_ _1156_
+ _1157_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__o22a_1
Xhold19 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] vssd1 vssd1 vccd1 vccd1 net476
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ clknet_leaf_18_wb_clk_i _0596_ _0124_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3043__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4056_ clknet_leaf_15_wb_clk_i _0541_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4663__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3007_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] net190 vssd1 vssd1 vccd1
+ vccd1 _1498_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout145_X net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4171__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3909_ net247 vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4140__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4290__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3189__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2240_ _1016_ _1017_ _1019_ _1021_ vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__or4b_1
XFILLER_0_57_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2171_ team_10_WB.instance_to_wrap.correct\[2\] team_10_WB.instance_to_wrap.gamelogic.rights\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3454__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1955_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] net147 vssd1 vssd1 vccd1
+ vccd1 _0876_ sky130_fd_sc_hd__or2_1
XANTENNA__4013__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1886_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 _0810_ sky130_fd_sc_hd__inv_2
X_4674_ net183 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2450__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4163__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3625_ net267 vssd1 vssd1 vccd1 vccd1 _0157_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3038__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_898 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3556_ net234 vssd1 vssd1 vccd1 vccd1 _0088_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2507_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1223_ vssd1 vssd1
+ vccd1 vccd1 _1224_ sky130_fd_sc_hd__or2_1
X_3487_ net241 vssd1 vssd1 vccd1 vccd1 _0019_ sky130_fd_sc_hd__inv_2
X_2438_ net720 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__a221o_1
X_2369_ _0871_ _1143_ _1087_ vssd1 vssd1 vccd1 vccd1 _1144_ sky130_fd_sc_hd__a21oi_1
X_4108_ clknet_leaf_10_wb_clk_i _0579_ _0107_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_4039_ clknet_leaf_21_wb_clk_i _0524_ _0080_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_746 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input35_A wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3436__B1 _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2239__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1998__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4036__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4186__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2270__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3410_ team_10_WB.instance_to_wrap.host_row1\[68\] _1703_ net180 team_10_WB.instance_to_wrap.host_row2\[60\]
+ _1785_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__a221o_1
X_4390_ clknet_leaf_5_wb_clk_i _0775_ _0373_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[27\]
+ sky130_fd_sc_hd__dfstp_1
X_3341_ team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] _1701_ net180 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\]
+ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__a22o_1
X_3272_ net297 _1661_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__nor2_1
X_2223_ net42 net40 net43 _1007_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__and4_1
X_2154_ _0822_ net218 _0948_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_37_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2085_ team_10_WB.instance_to_wrap.dispFSM.guesses\[27\] net113 net140 net723 vssd1
+ vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__o22a_1
XANTENNA__2445__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_wb_clk_i_X clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1989__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2987_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] net161 _1491_ net217
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[25\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_1027 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1938_ _0840_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__nand2_1
X_4657_ net426 vssd1 vssd1 vccd1 vccd1 la_data_out[27] sky130_fd_sc_hd__buf_2
X_1869_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] vssd1 vssd1 vccd1 vccd1
+ _0794_ sky130_fd_sc_hd__inv_2
XANTENNA__2953__A2 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3608_ net278 vssd1 vssd1 vccd1 vccd1 _0140_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4588_ net452 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XFILLER_0_12_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3539_ net233 vssd1 vssd1 vccd1 vccd1 _0071_ sky130_fd_sc_hd__inv_2
XANTENNA__4059__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4568__444 vssd1 vssd1 vccd1 vccd1 net444 _4568__444/LO sky130_fd_sc_hd__conb_1
XANTENNA__3418__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540__352 vssd1 vssd1 vccd1 vccd1 _4540__352/HI net352 sky130_fd_sc_hd__conb_1
XFILLER_0_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_X net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3409__B1 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2880__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2910_ net590 net156 net125 net599 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[15\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3890_ net277 vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__inv_2
X_2841_ _1010_ _1238_ _1241_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2772_ team_10_WB.instance_to_wrap.clock_div.count\[25\] team_10_WB.instance_to_wrap.clock_div.count\[24\]
+ team_10_WB.instance_to_wrap.clock_div.count\[26\] _1382_ vssd1 vssd1 vccd1 vccd1
+ _1386_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4511_ net323 vssd1 vssd1 vccd1 vccd1 ADR_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4442_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[39\]
+ _0425_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold116 team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] vssd1 vssd1 vccd1 vccd1
+ net573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold105 team_10_WB.instance_to_wrap.dispFSM.guesses\[13\] vssd1 vssd1 vccd1 vccd1
+ net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 team_10_WB.instance_to_wrap.host_row1\[69\] vssd1 vssd1 vccd1 vccd1 net584
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[7\] vssd1 vssd1 vccd1
+ vccd1 net606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 team_10_WB.instance_to_wrap.dispFSM.guesses\[79\] vssd1 vssd1 vccd1 vccd1
+ net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4373_ clknet_leaf_1_wb_clk_i _0758_ _0356_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3360__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _1681_ _1698_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__and2_2
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3255_ _0813_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4201__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2206_ net194 _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__nor2_2
XANTENNA__3840__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3186_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\]
+ _1608_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__and3_1
XANTENNA__3051__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2137_ net134 _0933_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2068_ team_10_WB.instance_to_wrap.dispFSM.guesses\[44\] net109 net135 net624 vssd1
+ vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__o22a_1
XANTENNA__4671__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4524__336 vssd1 vssd1 vccd1 vccd1 _4524__336/HI net336 sky130_fd_sc_hd__conb_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2926__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3351__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4611__386 vssd1 vssd1 vccd1 vccd1 _4611__386/HI net386 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_28_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4224__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3342__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output66_A net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3660__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4374__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] _1514_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[56\] sky130_fd_sc_hd__mux2_1
XFILLER_0_59_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3942_ net238 vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__inv_2
X_3873_ net267 vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__inv_2
X_2824_ _1418_ _1426_ _1407_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_822 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2908__A2 _1181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2755_ net732 _1374_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2686_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\]
+ _1332_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__and3_1
X_4425_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[22\]
+ _0408_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3333__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4356_ clknet_leaf_19_wb_clk_i _0746_ _0345_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_3307_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4666__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4287_ clknet_leaf_15_wb_clk_i _0677_ _0276_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3238_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ _1638_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout175_X net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3169_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1551_ _1595_ vssd1 vssd1 vccd1
+ vccd1 _0500_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_11_wb_clk_i_X clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4397__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3088__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_41_Left_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload14 clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__clkinv_2
Xclkload25 clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload25/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2540_ _0818_ _0842_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2471_ net568 net129 _1194_ _1209_ vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4210_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[72\]
+ _0199_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[72\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Left_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4141_ clknet_leaf_9_wb_clk_i _0612_ _0140_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_4072_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[3\]
+ _0092_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3023_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3925_ net248 vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3856_ net262 vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout135_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload8 clknet_leaf_30_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XFILLER_0_27_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2807_ _1413_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__inv_2
XANTENNA__3003__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3565__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3787_ net272 vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout302_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2738_ team_10_WB.instance_to_wrap.clock_div.count\[13\] team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ _1362_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__and3_1
X_4408_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[5\]
+ _0391_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2669_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] _1321_ _1319_ vssd1
+ vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__o21ai_1
Xfanout201 net63 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout223 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\] vssd1 vssd1 vccd1
+ vccd1 net223 sky130_fd_sc_hd__clkbuf_2
XANTENNA__4169__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout212 team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1
+ net212 sky130_fd_sc_hd__clkbuf_4
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_4
Xfanout245 net249 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_4
X_4339_ clknet_leaf_20_wb_clk_i _0729_ _0328_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[62\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout234 net239 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_4
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout289 net290 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__buf_4
Xfanout267 net283 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_4
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4412__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1971_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__o22a_1
X_3710_ net235 vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__inv_2
X_4690_ net438 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[29] sky130_fd_sc_hd__buf_2
X_3641_ net263 vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3572_ net264 vssd1 vssd1 vccd1 vccd1 _0104_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2744__B1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2523_ net530 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] vssd1 vssd1
+ vccd1 vccd1 _0522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2454_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] net186 vssd1 vssd1 vccd1
+ vccd1 _1200_ sky130_fd_sc_hd__or2_1
XANTENNA__1904__Y _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2385_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1157_ sky130_fd_sc_hd__a21o_1
X_4124_ clknet_leaf_17_wb_clk_i _0595_ _0123_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 gpio_in[24] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_4055_ clknet_leaf_15_wb_clk_i _0540_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_3006_ net212 net126 _1496_ net725 net158 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[39\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout252_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3908_ net264 vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3839_ net258 vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_641 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4435__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3189__B net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2170_ _0961_ _0960_ _0959_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_38_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3952__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4272__Q team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_1954_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4673_ net182 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4308__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1885_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 _0809_ sky130_fd_sc_hd__inv_2
X_3624_ net267 vssd1 vssd1 vccd1 vccd1 _0156_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2193__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3555_ net233 vssd1 vssd1 vccd1 vccd1 _0087_ sky130_fd_sc_hd__inv_2
X_3486_ _1409_ _1436_ _1438_ _1405_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__o211a_1
XANTENNA__3390__B1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2506_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2437_ net539 net132 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__a22o_1
XANTENNA__4458__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3054__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2368_ _1091_ _1137_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__xor2_1
X_4107_ clknet_leaf_2_wb_clk_i _0578_ _0106_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4674__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2299_ _1077_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__inv_2
XANTENNA__3445__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4038_ clknet_leaf_21_wb_clk_i _0523_ _0079_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2487__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3436__A1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2239__A2 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3975__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1998__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3340_ _1694_ _1718_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__nor2_4
XANTENNA__3663__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3372__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3271_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ vssd1 vssd1 vccd1 vccd1
+ _1661_ sky130_fd_sc_hd__and4_1
X_2222_ net182 vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__inv_2
XANTENNA__2478__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2153_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] net109 net136 net688 vssd1
+ vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4130__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2938__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2986_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] net164 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[24\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1937_ _0842_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3049__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4656_ net425 vssd1 vssd1 vccd1 vccd1 la_data_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_44_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1868_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1 vccd1 vccd1
+ _0793_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout215_A team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3607_ net261 vssd1 vssd1 vccd1 vccd1 _0139_ sky130_fd_sc_hd__inv_2
X_4587_ net200 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3573__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3538_ net233 vssd1 vssd1 vccd1 vccd1 _0070_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2189__A team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3469_ team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] net181 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[71\]
+ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__a22o_1
XANTENNA__2469__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3998__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_23_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2929__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3354__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_282 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4003__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3409__B2 team_10_WB.instance_to_wrap.host_row2\[84\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4153__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2840_ _1405_ _1426_ _1437_ _1410_ vssd1 vssd1 vccd1 vccd1 _0004_ sky130_fd_sc_hd__a211oi_1
XANTENNA__2562__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2771_ team_10_WB.instance_to_wrap.clock_div.count\[26\] _1384_ vssd1 vssd1 vccd1
+ vccd1 _1385_ sky130_fd_sc_hd__nor2_1
X_4510_ net322 vssd1 vssd1 vccd1 vccd1 ADR_O[17] sky130_fd_sc_hd__buf_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4441_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[38\]
+ _0424_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ sky130_fd_sc_hd__dfstp_1
Xhold106 _0680_ vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _0698_ vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\] vssd1 vssd1 vccd1
+ vccd1 net585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[4\] vssd1 vssd1 vccd1
+ vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4372_ clknet_leaf_6_wb_clk_i _0757_ _0355_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_3323_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ _1698_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__and3_4
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3254_ net706 _1609_ _1650_ net231 vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__o211a_1
X_2205_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] vssd1 vssd1 vccd1 vccd1 _0993_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3185_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\] vssd1 vssd1 vccd1 vccd1 _1608_
+ sky130_fd_sc_hd__and3_1
X_2136_ net217 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0933_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout165_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2067_ team_10_WB.instance_to_wrap.dispFSM.guesses\[53\] net143 net107 net565 vssd1
+ vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4563__375 vssd1 vssd1 vccd1 vccd1 _4563__375/HI net375 sky130_fd_sc_hd__conb_1
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2969_ net212 net126 _1482_ net689 net159 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[15\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2191__B team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout120_X net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4639_ net408 vssd1 vssd1 vccd1 vccd1 la_data_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__3336__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4026__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4176__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4547__359 vssd1 vssd1 vccd1 vccd1 _4547__359/HI net359 sky130_fd_sc_hd__conb_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3941_ net237 vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3872_ net268 vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__inv_2
X_2823_ _0514_ _0513_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2754_ _1373_ _1374_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[19\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4049__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2685_ _1334_ _1335_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[8\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4424_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[21\]
+ _0407_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4199__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4355_ clknet_leaf_19_wb_clk_i _0745_ _0344_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[78\]
+ sky130_fd_sc_hd__dfstp_1
X_3306_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_39_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4286_ clknet_leaf_17_wb_clk_i _0676_ _0275_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3062__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3237_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ _1637_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] vssd1 vssd1 vccd1 vccd1
+ _1641_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout282_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3168_ _1586_ _1590_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4682__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2119_ _0920_ _0921_ vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__nor2_1
X_3099_ _0789_ net207 vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout168_X net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3254__C1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_675 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_X clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4652__421 vssd1 vssd1 vccd1 vccd1 _4652__421/HI net421 sky130_fd_sc_hd__conb_1
XFILLER_0_25_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input10_A wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload26 clknet_leaf_13_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_12
Xclkload15 clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload15/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3012__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2470_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] net197 team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ _1191_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__a22o_1
X_4140_ clknet_leaf_9_wb_clk_i _0611_ _0139_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4491__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[2\]
+ _0091_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3022_ net501 net185 _1505_ net208 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[47\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__3484__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4275__Q team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_915 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2039__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3924_ net265 vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3855_ net277 vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload9 clknet_leaf_31_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__inv_16
X_2806_ net230 _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__nand2_1
X_3786_ net281 vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_2737_ team_10_WB.instance_to_wrap.clock_div.count\[13\] _1362_ net716 vssd1 vssd1
+ vccd1 vccd1 _1363_ sky130_fd_sc_hd__a21oi_1
X_4636__405 vssd1 vssd1 vccd1 vccd1 _4636__405/HI net405 sky130_fd_sc_hd__conb_1
X_2668_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] _1321_ vssd1 vssd1
+ vccd1 vccd1 _1324_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4407_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[4\]
+ _0390_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4677__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2599_ _0903_ _1280_ _1282_ vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__and3b_1
Xfanout213 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1 vccd1
+ net213 sky130_fd_sc_hd__clkbuf_4
Xfanout202 net209 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net249 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
Xfanout224 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] vssd1 vssd1 vccd1
+ vccd1 net224 sky130_fd_sc_hd__clkbuf_2
Xfanout235 net239 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_4
X_4338_ clknet_leaf_19_wb_clk_i net570 _0327_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[61\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout279 net283 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__buf_2
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__buf_4
XANTENNA_input2_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4269_ clknet_leaf_0_wb_clk_i _0659_ _0258_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4214__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4364__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_53_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1970_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] net150 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\]
+ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_23_Left_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2441__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2992__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3640_ net253 vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__inv_2
X_3571_ net271 vssd1 vssd1 vccd1 vccd1 _0103_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2522_ net496 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1
+ vccd1 vccd1 _0523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2453_ net601 net133 _1185_ _1199_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__a22o_1
X_2384_ _1154_ _1155_ _1087_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__a21oi_1
X_4123_ clknet_leaf_18_wb_clk_i _0594_ _0122_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_4054_ clknet_leaf_15_wb_clk_i _0539_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
X_3005_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\] net165 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[38\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3472__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4387__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout245_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3907_ net254 vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3838_ net259 vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2196__C1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3769_ net292 vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input5_X net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3463__A2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3311__A_N net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2974__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3151__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4665__431 vssd1 vssd1 vccd1 vccd1 _4665__431/HI net431 sky130_fd_sc_hd__conb_1
XANTENNA__3454__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1953_ net147 net157 vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4672_ net182 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2965__B2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1884_ team_10_WB.instance_to_wrap.message_reg.state\[0\] vssd1 vssd1 vccd1 vccd1
+ _0808_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3623_ net269 vssd1 vssd1 vccd1 vccd1 _0155_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3554_ net239 vssd1 vssd1 vccd1 vccd1 _0086_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_998 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3485_ net549 _1284_ _0885_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__o21a_1
X_2505_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1 _1222_
+ sky130_fd_sc_hd__and3b_1
X_2436_ _1193_ _1194_ net557 net132 vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2367_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] _1084_ _1140_
+ _1142_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__o22a_1
X_4106_ clknet_leaf_10_wb_clk_i _0577_ _0105_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2298_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _0823_ _1069_ vssd1 vssd1
+ vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand3_1
X_4037_ clknet_leaf_21_wb_clk_i _0522_ _0078_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3070__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3445__A2 _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout150_X net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_203 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3381__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4402__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A2 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4591__455 vssd1 vssd1 vccd1 vccd1 net455 _4591__455/LO sky130_fd_sc_hd__conb_1
X_3270_ net297 _1659_ _1660_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__nor3_1
X_2221_ _1001_ _1002_ _1003_ _1006_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__or4_1
X_2152_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__nor2_1
XANTENNA__2883__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2083_ net576 net143 net107 net607 vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1989__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2938__A1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2985_ _1491_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1936_ net229 _0857_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__or3b_2
XPHY_EDGE_ROW_26_Left_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4655_ net424 vssd1 vssd1 vccd1 vccd1 la_data_out[25] sky130_fd_sc_hd__buf_2
X_1867_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] vssd1 vssd1 vccd1 vccd1
+ _0792_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4425__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4586_ net200 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_1
X_3606_ net275 vssd1 vssd1 vccd1 vccd1 _0138_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout110_A net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout208_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3537_ net233 vssd1 vssd1 vccd1 vccd1 _0069_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_10_Left_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3065__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ net632 net177 _1841_ net230 vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__o211a_1
XANTENNA__2189__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3399_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] _1688_ _1679_ net210
+ vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__o211a_1
X_2419_ net202 _0942_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__and2_2
XANTENNA_fanout198_X net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2874__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2636__C _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3051__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input40_A wbs_cyc_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4368__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3409__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4448__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3042__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2770_ _1383_ _1384_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[25\]
+ sky130_fd_sc_hd__nor2_1
Xhold107 team_10_WB.instance_to_wrap.host_row1\[68\] vssd1 vssd1 vccd1 vccd1 net564
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4440_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[37\]
+ _0423_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold129 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[7\] vssd1 vssd1 vccd1
+ vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[2\] vssd1 vssd1 vccd1
+ vccd1 net575 sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ clknet_leaf_6_wb_clk_i _0756_ _0354_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3322_ _1683_ _1694_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nor2_1
X_3253_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] _1607_ _1609_ vssd1 vssd1
+ vccd1 vccd1 _1650_ sky130_fd_sc_hd__nand3_1
X_3184_ _1603_ _1604_ _1605_ _1606_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__or4_1
X_2204_ _0946_ net194 _0990_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__o21ai_1
X_2135_ net134 _0932_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__and2_1
X_2066_ team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] net111 net138 net637 vssd1
+ vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3849__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout158_A net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2472__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2968_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] net162 _1483_ net213
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[14\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1919_ team_10_WB.instance_to_wrap.host_col\[2\] team_10_WB.instance_to_wrap.host_col\[1\]
+ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__or3_2
X_4638_ net407 vssd1 vssd1 vccd1 vccd1 la_data_out[8] sky130_fd_sc_hd__buf_2
X_2899_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\] net155 net122 net612
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[4\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3965__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4569_ net445 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3024__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_28 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input43_X net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4120__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3940_ net265 vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3871_ net267 vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__inv_2
X_2822_ net282 _1417_ vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2753_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[19\]
+ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1367_ vssd1 vssd1 vccd1 vccd1
+ _1374_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2684_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1332_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4423_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[20\]
+ _0406_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_4354_ clknet_leaf_19_wb_clk_i _0744_ _0343_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_3305_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__and2b_2
X_4285_ clknet_leaf_14_wb_clk_i _0675_ _0274_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
X_3236_ net666 _1638_ _1640_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4530__342 vssd1 vssd1 vccd1 vccd1 _4530__342/HI net342 sky130_fd_sc_hd__conb_1
X_3167_ team_10_WB.instance_to_wrap.dispFSM.msg\[4\] _1278_ _1568_ _1593_ vssd1 vssd1
+ vccd1 vccd1 _1594_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3098_ net198 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] _0995_ _1543_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\] sky130_fd_sc_hd__o31a_1
X_2118_ team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] team_10_WB.instance_to_wrap.buffer.temp_guess\[6\]
+ team_10_WB.instance_to_wrap.buffer.temp_guess\[5\] team_10_WB.instance_to_wrap.buffer.temp_guess\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_1_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ net611 net145 net108 net645 vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_770 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_687 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4143__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3088__A3 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4293__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3489__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_662 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload16 clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload27 clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload27/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_24_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output71_A net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514__326 vssd1 vssd1 vccd1 vccd1 _4514__326/HI net326 sky130_fd_sc_hd__conb_1
XANTENNA__3016__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ clknet_leaf_22_wb_clk_i net491 _0090_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3021_ _0796_ net185 vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2039__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3923_ net248 vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__inv_2
X_3854_ net258 vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2805_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[1\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3785_ net292 vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__inv_2
XANTENNA__4166__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4675__433 vssd1 vssd1 vccd1 vccd1 _4675__433/HI net433 sky130_fd_sc_hd__conb_1
X_4601__376 vssd1 vssd1 vccd1 vccd1 _4601__376/HI net376 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_30_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2736_ net571 _1362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[13\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2667_ _1318_ _1322_ _1323_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[2\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_14_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1970__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4406_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[3\]
+ _0389_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout203 net209 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
X_2598_ _1275_ _1278_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__or2_1
Xfanout214 team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1 vccd1
+ net214 sky130_fd_sc_hd__buf_4
X_4337_ clknet_leaf_16_wb_clk_i _0727_ _0326_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[60\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 team_10_WB.instance_to_wrap.host_col\[2\] vssd1 vssd1 vccd1 vccd1 net225
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout236 net238 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_4
Xfanout247 net249 vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
Xfanout258 net260 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_4
X_4268_ clknet_leaf_3_wb_clk_i _0658_ _0257_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout269 net283 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_4
XANTENNA__2197__B net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\] _1628_ net172 vssd1
+ vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout180_X net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3475__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4199_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\]
+ _0188_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[61\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4039__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4189__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4659__428 vssd1 vssd1 vccd1 vccd1 _4659__428/HI net428 sky130_fd_sc_hd__conb_1
XANTENNA__2729__C1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3570_ net270 vssd1 vssd1 vccd1 vccd1 _0102_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2521_ net483 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] vssd1 vssd1
+ vccd1 vccd1 _0524_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1952__B1 _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2452_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] net186 vssd1 vssd1 vccd1
+ vccd1 _1199_ sky130_fd_sc_hd__or2_1
X_2383_ _1123_ _1127_ _1136_ _0871_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4122_ clknet_leaf_18_wb_clk_i _0593_ _0121_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_4053_ clknet_leaf_14_wb_clk_i _0538_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3004_ _1484_ _1496_ _1497_ _1493_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[37\]
+ sky130_fd_sc_hd__a22oi_1
Xinput3 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3906_ net259 vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout238_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3068__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_930 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2480__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3837_ net248 vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3768_ net293 vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__inv_2
X_2719_ _1351_ _1352_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__4688__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3699_ net236 vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3448__B1 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4481__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3384__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3007__A team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3439__A0 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2111__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1952_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0874_ _0873_ _0863_ vssd1
+ vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4671_ net182 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1883_ team_10_WB.instance_to_wrap.message_reg.state\[1\] vssd1 vssd1 vccd1 vccd1
+ _0807_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3622_ net269 vssd1 vssd1 vccd1 vccd1 _0154_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3553_ net289 vssd1 vssd1 vccd1 vccd1 _0085_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3484_ net71 net177 _1856_ net230 vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2504_ net223 _1221_ _1217_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__mux2_1
XANTENNA__4204__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2435_ net132 _1190_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4105_ clknet_leaf_8_wb_clk_i _0576_ _0104_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_2366_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout188_A net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2297_ _1069_ _1074_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__or2_1
XANTENNA__4354__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4036_ clknet_leaf_21_wb_clk_i _0521_ _0077_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_56_Left_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2653__B2 _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4607__382 vssd1 vssd1 vccd1 vccd1 _4607__382/HI net382 sky130_fd_sc_hd__conb_1
XANTENNA_30 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3497__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3372__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4377__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2220_ net32 net31 _1004_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__or4_1
X_2151_ net166 _0918_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__or2_1
X_2082_ team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] net111 net139 net669 vssd1
+ vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_37_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2984_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] net126 _1489_ _1490_
+ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__nand4_4
XFILLER_0_8_437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1935_ _0847_ net196 vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__nand2_2
XFILLER_0_12_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4654_ net423 vssd1 vssd1 vccd1 vccd1 la_data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_47_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1866_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] vssd1 vssd1 vccd1 vccd1
+ _0791_ sky130_fd_sc_hd__inv_2
X_3605_ net278 vssd1 vssd1 vccd1 vccd1 _0137_ sky130_fd_sc_hd__inv_2
X_4585_ net200 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3536_ net233 vssd1 vssd1 vccd1 vccd1 _0068_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3467_ net169 _1839_ _1840_ _1838_ _1403_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3398_ team_10_WB.instance_to_wrap.host_row2\[43\] team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__mux2_1
X_2418_ _1178_ _1179_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2349_ _1122_ _1102_ _1117_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__and3b_1
XANTENNA__3081__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4019_ clknet_leaf_28_wb_clk_i _0504_ _0066_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.unlocked
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3354__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input33_A wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 team_10_WB.instance_to_wrap.dispFSM.guesses\[45\] vssd1 vssd1 vccd1 vccd1
+ net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold119 team_10_WB.instance_to_wrap.dispFSM.guesses\[37\] vssd1 vssd1 vccd1 vccd1
+ net576 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ clknet_leaf_26_wb_clk_i _0755_ _0353_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3321_ _1686_ _1695_ vssd1 vssd1 vccd1 vccd1 _1701_ sky130_fd_sc_hd__and2_2
XFILLER_0_42_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3252_ _1610_ _1649_ net296 vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3183_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[12\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__or4bb_1
X_2203_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.correct\[0\]
+ team_10_WB.instance_to_wrap.correct\[2\] vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__and3b_2
XANTENNA__1922__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2134_ net216 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0932_ sky130_fd_sc_hd__mux2_1
X_2065_ team_10_WB.instance_to_wrap.dispFSM.guesses\[55\] net144 net107 net558 vssd1
+ vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ _1479_ _1483_ _1484_ _1482_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[13\]
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_60_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2898_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\] net155 net122 net609
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[3\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1918_ team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__nand2b_2
X_4637_ net406 vssd1 vssd1 vccd1 vccd1 la_data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_60_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3336__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3076__S net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4568_ net444 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
X_4499_ net311 vssd1 vssd1 vccd1 vccd1 ADR_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ net245 vssd1 vssd1 vccd1 vccd1 _0051_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4072__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4415__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4627__396 vssd1 vssd1 vccd1 vccd1 _4627__396/HI net396 sky130_fd_sc_hd__conb_1
XFILLER_0_14_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3870_ net267 vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__inv_2
X_2821_ _1405_ _1424_ _1425_ _1411_ _1419_ vssd1 vssd1 vccd1 vccd1 _0000_ sky130_fd_sc_hd__a32o_1
XANTENNA__3685__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2752_ net729 _1372_ vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2683_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[8\] _1332_ vssd1 vssd1
+ vccd1 vccd1 _1334_ sky130_fd_sc_hd__and2_1
X_4422_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[19\]
+ _0405_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4353_ clknet_leaf_16_wb_clk_i _0743_ _0342_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[76\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3304_ _0815_ net211 _1679_ _1681_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4284_ clknet_leaf_19_wb_clk_i net509 _0273_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3235_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\] _1638_ net172 vssd1
+ vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4095__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _0891_ _0899_ _0906_ net228 vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__and4bb_1
X_3097_ team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] net202 vssd1 vssd1 vccd1
+ vccd1 _1543_ sky130_fd_sc_hd__or2_1
X_2117_ team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] team_10_WB.instance_to_wrap.buffer.temp_guess\[2\]
+ team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] team_10_WB.instance_to_wrap.buffer.temp_guess\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__or4_1
X_2048_ team_10_WB.instance_to_wrap.dispFSM.guesses\[64\] net113 net140 net684 vssd1
+ vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3006__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3999_ clknet_leaf_25_wb_clk_i net458 net271 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2004__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4438__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload17 clknet_leaf_20_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_12
XFILLER_0_50_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload28 clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4553__365 vssd1 vssd1 vccd1 vccd1 _4553__365/HI net365 sky130_fd_sc_hd__conb_1
XANTENNA__3484__A1 net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3020_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[6\] net185 _1504_ net206
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[46\] sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3955__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3922_ net242 vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3853_ net238 vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__inv_2
X_2804_ _1405_ _1410_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3784_ net293 vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__inv_2
X_2735_ _1361_ _1362_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2666_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1323_ sky130_fd_sc_hd__a21o_1
XANTENNA__1970__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1970__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4405_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[2\]
+ _0388_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout204 net209 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_4
X_4336_ clknet_leaf_16_wb_clk_i _0726_ _0325_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[59\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2597_ _1275_ _1278_ vssd1 vssd1 vccd1 vccd1 _1282_ sky130_fd_sc_hd__nor2_1
Xfanout226 team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1 net226
+ sky130_fd_sc_hd__clkbuf_2
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_4
Xfanout215 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1 vccd1
+ net215 sky130_fd_sc_hd__buf_4
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__buf_4
X_4267_ clknet_leaf_4_wb_clk_i _0657_ _0256_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1950__X _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 net249 vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_4
X_4198_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[60\]
+ _0187_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[60\] sky130_fd_sc_hd__dfrtp_1
X_3218_ net713 _1626_ _1629_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_31_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_3149_ _0903_ _1277_ _1280_ _1578_ vssd1 vssd1 vccd1 vccd1 _1579_ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout173_X net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4110__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4496__308 vssd1 vssd1 vccd1 vccd1 _4496__308/HI net308 sky130_fd_sc_hd__conb_1
XFILLER_0_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4537__349 vssd1 vssd1 vccd1 vccd1 _4537__349/HI net349 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_53_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2910__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3978__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4392__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2441__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3439__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2520_ net524 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1
+ vccd1 vccd1 _0525_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2451_ net593 net131 _1185_ _1198_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2382_ _1123_ _1136_ _1127_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2901__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4121_ clknet_leaf_26_wb_clk_i _0592_ _0120_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_X clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4052_ clknet_leaf_15_wb_clk_i _0537_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_3003_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\] net161 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[4\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[36\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_2
XFILLER_0_36_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4133__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4642__411 vssd1 vssd1 vccd1 vccd1 _4642__411/HI net411 sky130_fd_sc_hd__conb_1
X_3905_ net257 vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3836_ net264 vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3767_ net280 vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__inv_2
XANTENNA__4283__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3393__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2718_ team_10_WB.instance_to_wrap.clock_div.count\[6\] _1349_ vssd1 vssd1 vccd1
+ vccd1 _1352_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3698_ net236 vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3084__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2649_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4319_ clknet_leaf_16_wb_clk_i _0709_ _0308_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_972 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3007__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1951_ team_10_WB.instance_to_wrap.host_message_reg.Cstate team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] _0861_ vssd1 vssd1 vccd1 vccd1
+ _0874_ sky130_fd_sc_hd__nor4_4
X_4670_ net184 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_1
X_1882_ team_10_WB.EN_VAL_REG vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
XFILLER_0_43_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3621_ net251 vssd1 vssd1 vccd1 vccd1 _0153_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3375__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3552_ net289 vssd1 vssd1 vccd1 vccd1 _0084_ sky130_fd_sc_hd__inv_2
XANTENNA__3693__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1925__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2503_ net223 _0889_ net222 vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__and3b_1
XFILLER_0_12_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4559__371 vssd1 vssd1 vccd1 vccd1 _4559__371/HI net371 sky130_fd_sc_hd__conb_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3483_ _1847_ _1853_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2434_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] _1192_ vssd1 vssd1 vccd1
+ vccd1 _1193_ sky130_fd_sc_hd__nor2_1
X_2365_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _0823_ _1069_ _1085_
+ vssd1 vssd1 vccd1 vccd1 _1141_ sky130_fd_sc_hd__a31o_1
X_4104_ clknet_leaf_25_wb_clk_i _0575_ _0103_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2296_ _0841_ _1069_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__or2_2
X_4035_ clknet_leaf_21_wb_clk_i _0520_ _0076_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3079__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_31 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3819_ net253 vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__inv_2
XANTENNA__3366__B1 _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4029__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout303_X net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2012__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4179__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3778__A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3357__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3018__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2150_ net166 _0918_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nor2_1
X_2081_ team_10_WB.instance_to_wrap.dispFSM.guesses\[39\] net144 net108 net573 vssd1
+ vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2983_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[24\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\]
+ _0836_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net160 vssd1 vssd1 vccd1
+ vccd1 _1490_ sky130_fd_sc_hd__a41o_1
XFILLER_0_9_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1934_ _0843_ net196 vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4653_ net422 vssd1 vssd1 vccd1 vccd1 la_data_out[23] sky130_fd_sc_hd__buf_2
Xinput40 wbs_cyc_i vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_1
X_1865_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] vssd1 vssd1 vccd1 vccd1
+ _0790_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2531__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3604_ net263 vssd1 vssd1 vccd1 vccd1 _0136_ sky130_fd_sc_hd__inv_2
X_4584_ net200 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_742 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3535_ net233 vssd1 vssd1 vccd1 vccd1 _0067_ sky130_fd_sc_hd__inv_2
XANTENNA__4321__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3466_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _1686_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ net210 vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__and4b_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2417_ _1164_ _1167_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout298_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3397_ team_10_WB.instance_to_wrap.host_row1\[59\] net169 _1768_ _1773_ vssd1 vssd1
+ vccd1 vccd1 _1774_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2348_ _1102_ _1117_ _1122_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__and3b_1
X_2279_ _0917_ _0948_ _1034_ _1047_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__o31ai_1
X_4018_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[2\]
+ net288 vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_419 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4344__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 _0712_ vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ team_10_WB.instance_to_wrap.host_row2\[40\] net174 _1699_ team_10_WB.instance_to_wrap.host_row1\[48\]
+ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3251_ _1609_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__nand2b_1
X_3182_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] vssd1 vssd1 vccd1 vccd1 _1605_
+ sky130_fd_sc_hd__or3b_1
X_2202_ _0918_ _0972_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2133_ net134 _0931_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__and2_1
X_2064_ team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] net113 net140 net711 vssd1
+ vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] _1192_ vssd1 vssd1 vccd1
+ vccd1 _1484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2897_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\] net153 net121 net604
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[2\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1917_ team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__and2b_1
X_4636_ net405 vssd1 vssd1 vccd1 vccd1 la_data_out[6] sky130_fd_sc_hd__buf_2
XFILLER_0_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout213_A team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4567_ net443 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
XFILLER_0_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4498_ net310 vssd1 vssd1 vccd1 vccd1 ADR_O[5] sky130_fd_sc_hd__buf_2
X_3518_ net246 vssd1 vssd1 vccd1 vccd1 _0050_ sky130_fd_sc_hd__inv_2
X_3449_ _1821_ _1822_ _1823_ net304 vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__o31a_1
XFILLER_0_58_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4217__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2960__A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4367__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3015__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2820_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2751_ _1371_ _1372_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[18\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2682_ _1318_ _1331_ _1333_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[7\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_5_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_901 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4421_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[18\]
+ _0404_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4352_ clknet_leaf_17_wb_clk_i _0742_ _0341_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[75\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2526__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3303_ _1680_ _1683_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__nor2_1
X_4283_ clknet_leaf_19_wb_clk_i _0673_ _0272_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3234_ net537 _1637_ _1639_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__o21a_1
X_3165_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1551_ _1591_ _1592_ vssd1 vssd1
+ vccd1 vccd1 _0499_ sky130_fd_sc_hd__o22a_1
X_3096_ net204 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[44\] net187 _1542_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[84\] sky130_fd_sc_hd__a31o_1
X_2116_ net157 _0918_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__or2_1
X_2047_ team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] net110 net137 net712 vssd1
+ vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3006__A2 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3998_ clknet_leaf_25_wb_clk_i net460 net271 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
X_2949_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] net162 _1478_ net217 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[1\] sky130_fd_sc_hd__o22a_1
XFILLER_0_44_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1973__C1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout216_X net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4619_ net391 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4007__RESET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2453__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload29 clknet_leaf_16_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__inv_6
Xclkload18 clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload18/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3484__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3313__X _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4564__440 vssd1 vssd1 vccd1 vccd1 net440 _4564__440/LO sky130_fd_sc_hd__conb_1
XFILLER_0_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3921_ net242 vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__inv_2
XANTENNA__2444__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3852_ net259 vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2803_ _1407_ _0517_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3783_ net281 vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2734_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] _1356_ vssd1 vssd1 vccd1 vccd1
+ _1362_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2665_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__inv_2
XANTENNA__1970__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4404_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[1\]
+ _0387_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_2596_ _1276_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand2_1
Xfanout205 net209 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
XANTENNA__4062__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4335_ clknet_leaf_15_wb_clk_i _0725_ _0324_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[58\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout238 net239 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_2
Xfanout227 _0897_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__clkbuf_2
Xfanout216 team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1 vccd1
+ net216 sky130_fd_sc_hd__buf_4
X_4266_ clknet_leaf_4_wb_clk_i _0656_ _0255_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout249 net266 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
X_3217_ net172 _1628_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__nor2_1
X_4197_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[59\]
+ _0186_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[59\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout280_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3475__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3148_ _1571_ _1577_ _1560_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3350__C_N net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3079_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout166_X net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2986__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4405__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 team_10_WB.instance_to_wrap.dispFSM.guesses\[24\] vssd1 vssd1 vccd1 vccd1
+ net727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2977__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4520__332 vssd1 vssd1 vccd1 vccd1 _4520__332/HI net332 sky130_fd_sc_hd__conb_1
XANTENNA__4085__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2450_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[26\] net185 vssd1 vssd1 vccd1
+ vccd1 _1198_ sky130_fd_sc_hd__or2_1
XANTENNA__1952__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2381_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] _1084_ _1141_
+ _1153_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__o22a_1
X_4120_ clknet_leaf_2_wb_clk_i _0591_ _0119_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_4051_ clknet_leaf_15_wb_clk_i _0536_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3457__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3002_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\] net162 _1497_ net215
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[35\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput5 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_2
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_6_wb_clk_i_X clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2968__B2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3904_ net257 vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1939__A team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2534__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4428__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ net247 vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3766_ net296 vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout126_A _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3393__A1 team_10_WB.instance_to_wrap.host_row2\[83\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2717_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ team_10_WB.instance_to_wrap.clock_div.count\[6\] _1347_ vssd1 vssd1 vccd1 vccd1
+ _1351_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3365__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3697_ net234 vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2648_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] team_10_WB.instance_to_wrap.uart_receiver.state\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.state\[1\] vssd1 vssd1 vccd1 vccd1 _1310_
+ sky130_fd_sc_hd__or3b_2
X_2579_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[1\] _1259_ _0904_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__o2bb2a_1
X_4318_ clknet_leaf_17_wb_clk_i _0708_ _0307_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4249_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[5\]
+ _0238_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3448__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3081__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4504__316 vssd1 vssd1 vccd1 vccd1 _4504__316/HI net316 sky130_fd_sc_hd__conb_1
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3384__A1 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_19 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3945__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2895__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_X net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2207__X _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1950_ _0841_ _0871_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__or2_2
XFILLER_0_56_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1881_ team_10_WB.instance_to_wrap.gamelogic.green vssd1 vssd1 vccd1 vccd1 _0806_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3620_ net269 vssd1 vssd1 vccd1 vccd1 _0152_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3551_ net289 vssd1 vssd1 vccd1 vccd1 _0083_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2502_ net626 _1220_ _1217_ vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3482_ _1727_ _1854_ _1403_ _1689_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2433_ net561 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2364_ _1138_ _1139_ _1088_ vssd1 vssd1 vccd1 vccd1 _1140_ sky130_fd_sc_hd__o21a_1
X_4103_ clknet_leaf_25_wb_clk_i _0574_ _0102_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__2529__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4100__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2295_ _0840_ _1073_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__nand2_2
XFILLER_0_56_1120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4034_ clknet_leaf_21_wb_clk_i _0519_ _0075_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.message_reg.msg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout243_A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3818_ net247 vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__inv_2
XANTENNA__3968__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_X net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3749_ net285 vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2012__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2877__A0 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4649__418 vssd1 vssd1 vccd1 vccd1 _4649__418/HI net418 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_39_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2644__A3 _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3357__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4123__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2080_ team_10_WB.instance_to_wrap.dispFSM.guesses\[32\] net113 net140 team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3321__X _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2979__A1_N _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2982_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[25\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] _0837_ net161 vssd1 vssd1 vccd1
+ vccd1 _1489_ sky130_fd_sc_hd__a41o_1
XFILLER_0_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1933_ _0850_ net196 vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4652_ net421 vssd1 vssd1 vccd1 vccd1 la_data_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__2812__S net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput30 wbs_adr_i[2] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_1
X_1864_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1 vccd1 vccd1
+ _0789_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3603_ net262 vssd1 vssd1 vccd1 vccd1 _0135_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4583_ net451 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
Xinput41 wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_656 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_678 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3534_ net251 vssd1 vssd1 vccd1 vccd1 _0066_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3465_ team_10_WB.instance_to_wrap.host_row1\[62\] team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload28_A clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2416_ _1177_ net232 _0849_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__and3b_2
X_3396_ team_10_WB.instance_to_wrap.host_row1\[43\] _1693_ _1770_ _1771_ _1772_ vssd1
+ vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__a2111o_1
X_2347_ _1117_ _1122_ vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__nand2_1
X_2278_ _0950_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__nor2_1
X_4017_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[1\]
+ net288 vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3036__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4146__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4620__392 vssd1 vssd1 vccd1 vccd1 _4620__392/HI net392 sky130_fd_sc_hd__conb_1
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input19_A wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_507 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2250__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3250_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\] _1608_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__a21o_1
X_3181_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[19\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[18\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\]
+ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__or4b_1
XFILLER_0_28_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2201_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] _0989_ _0973_ vssd1
+ vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o21a_1
X_2132_ net215 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2063_ team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] net109 net135 net683 vssd1
+ vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__o22a_1
XANTENNA__4019__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2965_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\] net163 _1483_ net214
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[12\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__1947__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2542__S _1179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4169__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2896_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\] net154 net122 net619
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[1\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1916_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ _0839_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ net404 vssd1 vssd1 vccd1 vccd1 la_data_out[5] sky130_fd_sc_hd__buf_2
X_4566_ net442 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XANTENNA_fanout206_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3517_ net245 vssd1 vssd1 vccd1 vccd1 _0049_ sky130_fd_sc_hd__inv_2
X_4497_ net309 vssd1 vssd1 vccd1 vccd1 ADR_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3448_ team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] net171 _1704_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1823_ sky130_fd_sc_hd__a22o_1
X_3379_ team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] net173 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[2\]
+ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__a221o_1
X_4685__437 vssd1 vssd1 vccd1 vccd1 _4685__437/HI net437 sky130_fd_sc_hd__conb_1
XFILLER_0_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_3__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_62_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_781 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1991__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2215__X _1001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2750_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1365_ vssd1 vssd1 vccd1 vccd1
+ _1372_ sky130_fd_sc_hd__and4_1
XANTENNA__4461__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2681_ _1332_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4420_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[17\]
+ _0403_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4351_ clknet_leaf_16_wb_clk_i _0741_ _0340_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[74\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3302_ _1681_ _1682_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__nand2_1
X_4282_ clknet_leaf_18_wb_clk_i net485 _0271_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3233_ net172 _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__nor2_1
X_3164_ team_10_WB.instance_to_wrap.dispFSM.msg\[3\] _1278_ _1568_ _0903_ vssd1 vssd1
+ vccd1 vccd1 _1592_ sky130_fd_sc_hd__a211o_1
X_3095_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] net198 vssd1 vssd1 vccd1
+ vccd1 _1542_ sky130_fd_sc_hd__and2_1
X_2115_ _0916_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__or2_2
X_2046_ team_10_WB.instance_to_wrap.dispFSM.guesses\[66\] net111 net138 net640 vssd1
+ vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout156_A _1181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3997_ clknet_leaf_24_wb_clk_i _0487_ _0065_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2948_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] net165 _1478_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[0\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_356 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4618_ net390 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XANTENNA__3892__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2879_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net224 vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__and3b_1
XANTENNA__2517__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_X net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4549_ net361 vssd1 vssd1 vccd1 vccd1 DAT_O[23] sky130_fd_sc_hd__buf_2
XFILLER_0_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3478__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4334__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4484__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1964__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload19 clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_2_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3469__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3920_ net240 vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3851_ net248 vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__inv_2
X_2802_ _1409_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__inv_2
X_3782_ net295 vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__inv_2
X_2733_ team_10_WB.instance_to_wrap.clock_div.count\[12\] _1360_ vssd1 vssd1 vccd1
+ vccd1 _1361_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2664_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\] vssd1 vssd1 vccd1 vccd1
+ _1321_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4207__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4403_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[0\]
+ _0386_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2595_ _0908_ _1279_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4334_ clknet_leaf_17_wb_clk_i _0724_ _0323_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[57\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout206 net208 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
Xfanout228 _0897_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout217 team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1 vccd1
+ net217 sky130_fd_sc_hd__buf_4
XANTENNA__4357__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4265_ clknet_leaf_4_wb_clk_i _0655_ _0254_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload10_A clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout239 net266 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
X_3216_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] _1626_ vssd1 vssd1 vccd1
+ vccd1 _1628_ sky130_fd_sc_hd__and2_1
X_4196_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[58\]
+ _0185_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[58\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2132__A0 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3147_ _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout273_A net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ team_10_WB.instance_to_wrap.gamelogic.setWord\[27\] _1533_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[75\] sky130_fd_sc_hd__mux2_1
X_2029_ net195 _0909_ _0911_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout159_X net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_17_Left_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold260 net64 vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] vssd1 vssd1 vccd1 vccd1
+ net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2910__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2966__A team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2380_ _0871_ _1088_ _1152_ _1075_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__a32o_1
XANTENNA__2901__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3324__X _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ clknet_leaf_14_wb_clk_i _0535_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_3001_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\] net162 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[2\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[34\]
+ sky130_fd_sc_hd__o22a_1
Xinput6 gpio_in[37] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_1
XFILLER_0_36_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ net278 vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3834_ net259 vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2116__A net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3765_ net285 vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1955__A team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3393__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2716_ _1171_ _1349_ _1350_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[5\]
+ sky130_fd_sc_hd__nor3_1
X_3696_ net234 vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2647_ _1307_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2578_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] _0898_ _0901_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4317_ clknet_leaf_12_wb_clk_i _0707_ _0306_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[40\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3381__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4248_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[4\]
+ _0237_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4179_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[41\]
+ _0168_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[41\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4543__355 vssd1 vssd1 vccd1 vccd1 _4543__355/HI net355 sky130_fd_sc_hd__conb_1
XFILLER_0_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4014__Q team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3384__A2 net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_502 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4052__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1880_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1 vccd1
+ _0805_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3319__X _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3375__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ net286 vssd1 vssd1 vccd1 vccd1 _0082_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2501_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3481_ team_10_WB.instance_to_wrap.host_row2\[71\] team_10_WB.instance_to_wrap.dispFSM.guesses\[47\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2432_ net194 _1186_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__or2_1
X_2363_ net229 _0847_ _0853_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__and3b_1
XANTENNA__2886__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4102_ clknet_leaf_25_wb_clk_i _0573_ _0101_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4033_ clknet_leaf_10_wb_clk_i _0518_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_2294_ _0859_ _0865_ _1071_ _1072_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1007 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4527__339 vssd1 vssd1 vccd1 vccd1 _4527__339/HI net339 sky130_fd_sc_hd__conb_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_760 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ net256 vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3748_ net286 vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3679_ net242 vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3108__C net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4075__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4009__Q team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3357__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4632__401 vssd1 vssd1 vccd1 vccd1 _4632__401/HI net401 sky130_fd_sc_hd__conb_1
XANTENNA__4418__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ net212 _1485_ _1488_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[23\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1932_ team_10_WB.instance_to_wrap.host_col\[3\] net225 net226 team_10_WB.instance_to_wrap.host_col\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4651_ net420 vssd1 vssd1 vccd1 vccd1 la_data_out[21] sky130_fd_sc_hd__buf_2
XFILLER_0_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1863_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] vssd1 vssd1 vccd1 vccd1
+ _0788_ sky130_fd_sc_hd__inv_2
X_3602_ net276 vssd1 vssd1 vccd1 vccd1 _0134_ sky130_fd_sc_hd__inv_2
Xinput20 wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput31 wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_4582_ net450 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
Xinput42 wbs_stb_i vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_4
XFILLER_0_4_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3533_ net270 vssd1 vssd1 vccd1 vccd1 _0065_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3464_ _1828_ _1831_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2415_ net232 _1171_ net459 vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3395_ team_10_WB.instance_to_wrap.host_row1\[51\] _1699_ net179 team_10_WB.instance_to_wrap.host_row2\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4098__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2346_ _0829_ _1121_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\] vssd1 vssd1
+ vccd1 vccd1 _1122_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout186_A _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2277_ _1054_ _1055_ _1058_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__and3b_1
X_4016_ clknet_leaf_23_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[0\]
+ net288 vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_2__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_2__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4206__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4549__361 vssd1 vssd1 vccd1 vccd1 _4549__361/HI net361 sky130_fd_sc_hd__conb_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2200_ net134 _0971_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a21oi_1
X_3180_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\]
+ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__or4b_1
X_2131_ net134 _0930_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2062_ team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] net111 net141 net714 vssd1
+ vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__o22a_1
XANTENNA__3958__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2964_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] net161 _1483_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[11\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1915_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] vssd1 vssd1 vccd1 vccd1
+ _0838_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4678__434 vssd1 vssd1 vccd1 vccd1 _4678__434/HI net434 sky130_fd_sc_hd__conb_1
X_2895_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\] net155 net122 net622
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[0\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4634_ net403 vssd1 vssd1 vccd1 vccd1 la_data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_0_44_368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4565_ net441 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3516_ net245 vssd1 vssd1 vccd1 vccd1 _0048_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4496_ net308 vssd1 vssd1 vccd1 vccd1 ADR_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3447_ team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] net175 net168 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\]
+ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a22o_1
X_3378_ team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] _1715_ _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[66\]
+ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2329_ _0819_ _0849_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[1\] vssd1
+ vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout189_X net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2018__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4113__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1991__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1873__A team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2940__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_31_Left_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input31_A wbs_adr_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2456__C1 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2471__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2680_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\]
+ _1327_ vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4350_ clknet_leaf_17_wb_clk_i _0740_ _0339_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[73\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3301_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net211 vssd1 vssd1 vccd1
+ vccd1 _1682_ sky130_fd_sc_hd__nor2_1
XANTENNA__2931__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4281_ clknet_leaf_14_wb_clk_i _0671_ _0270_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3232_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] _1637_ vssd1 vssd1 vccd1
+ vccd1 _1638_ sky130_fd_sc_hd__and2_1
X_3163_ _1586_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__xor2_1
X_2114_ net219 net218 vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__nand2_1
X_3094_ net204 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] net187 _1541_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[83\] sky130_fd_sc_hd__a31o_1
X_2045_ team_10_WB.instance_to_wrap.dispFSM.guesses\[67\] net110 net137 team_10_WB.instance_to_wrap.dispFSM.guesses\[75\]
+ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__o22a_1
XANTENNA__4136__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2462__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3996_ clknet_leaf_24_wb_clk_i _0486_ _0064_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2947_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[1\] net165 _1475_ _1476_ _1477_
+ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_44_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4286__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3946__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4617_ net389 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2878_ net193 _1462_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[2\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4548_ net360 vssd1 vssd1 vccd1 vccd1 DAT_O[22] sky130_fd_sc_hd__buf_2
XFILLER_0_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4479_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[36\]
+ _0462_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2922__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_382 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1868__A team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4016__RESET_B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1964__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1964__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4009__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2913__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4159__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3850_ net242 vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2801_ net231 _1408_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3781_ net272 vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2732_ _1359_ _1360_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[11\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2663_ net533 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\] _1320_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2594_ _0890_ net228 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\] vssd1
+ vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4402_ clknet_leaf_1_wb_clk_i _0787_ _0385_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[39\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__2904__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4333_ clknet_leaf_14_wb_clk_i _0723_ _0322_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[56\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__buf_2
X_4264_ clknet_leaf_4_wb_clk_i _0654_ _0253_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout218 team_10_WB.instance_to_wrap.gamelogic.state\[1\] vssd1 vssd1 vccd1 vccd1
+ net218 sky130_fd_sc_hd__buf_2
Xfanout229 _0846_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_2
XANTENNA__2380__B2 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3215_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\] _1624_ _1627_ _1611_
+ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4195_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[57\]
+ _0184_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[57\] sky130_fd_sc_hd__dfrtp_1
X_3146_ _1573_ _1574_ _1569_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__a21oi_1
X_3077_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout266_A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2028_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3396__B1 _1770_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[16\]
+ _0047_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold261 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1
+ net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 team_10_WB.instance_to_wrap.clock_div.count\[25\] vssd1 vssd1 vccd1 vccd1
+ net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4301__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold272 team_10_WB.instance_to_wrap.clock_div.count\[19\] vssd1 vssd1 vccd1 vccd1
+ net729 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2371__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__B1 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4451__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2206__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3387__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2222__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3000_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\] net161 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[1\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[33\]
+ sky130_fd_sc_hd__o22a_1
Xinput7 wb_rst_i vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3902_ net259 vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3833_ net257 vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3378__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3764_ net291 vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2715_ team_10_WB.instance_to_wrap.clock_div.count\[4\] _1347_ team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__a21oi_1
X_3695_ net233 vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__inv_2
XANTENNA__1955__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2646_ team_10_WB.instance_to_wrap.uart_receiver.state\[2\] _0827_ team_10_WB.instance_to_wrap.uart_receiver.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__or3_1
XANTENNA__4324__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2577_ _1254_ _1255_ _1260_ _1261_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__o211a_1
X_4316_ clknet_leaf_18_wb_clk_i _0706_ _0305_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4474__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4247_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[3\]
+ _0236_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4178_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[40\]
+ _0167_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[40\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4209__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3129_ _1557_ _1559_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2895__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4205__Q team_10_WB.instance_to_wrap.host_row2\[67\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4347__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2500_ net220 net222 net223 net221 vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__or4b_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3480_ team_10_WB.instance_to_wrap.host_row2\[55\] net170 _1848_ _1852_ vssd1 vssd1
+ vccd1 vccd1 _1853_ sky130_fd_sc_hd__a211o_1
X_2431_ net194 _1186_ vssd1 vssd1 vccd1 vccd1 _1191_ sky130_fd_sc_hd__nor2_2
XFILLER_0_11_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2362_ _1091_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2293_ _0843_ net229 net196 _0858_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__nand4b_1
X_4101_ clknet_leaf_24_wb_clk_i _0572_ _0100_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4032_ clknet_leaf_12_wb_clk_i _0517_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_1__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3070__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_12 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2414__X _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_772 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3816_ net247 vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3747_ net272 vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ net240 vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2629_ _0807_ _0808_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.blue sky130_fd_sc_hd__nor2_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4510__322 vssd1 vssd1 vccd1 vccd1 _4510__322/HI net322 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_39_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1876__A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2980_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[22\] net160 _1488_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[22\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1931_ net229 _0848_ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1
+ vccd1 _0854_ sky130_fd_sc_hd__o21a_1
X_4650_ net419 vssd1 vssd1 vccd1 vccd1 la_data_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_51_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 wbs_adr_i[11] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_3601_ net276 vssd1 vssd1 vccd1 vccd1 _0133_ sky130_fd_sc_hd__inv_2
Xinput21 wbs_adr_i[21] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
Xinput43 wbs_we_i vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_4
X_4581_ net199 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput32 wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3532_ net270 vssd1 vssd1 vccd1 vccd1 _0064_ sky130_fd_sc_hd__inv_2
X_3463_ team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] net179 _1832_ _1836_ vssd1
+ vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__a211o_1
XANTENNA__2308__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2414_ team_10_WB.instance_to_wrap.clock_div.count\[6\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ _1170_ _1176_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__or4_4
XFILLER_0_0_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3394_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net210 _1681_ _1686_
+ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2345_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _0870_ _1118_ _1120_
+ _0828_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__a32o_1
X_2276_ _0791_ net212 _1050_ _1053_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__o2111a_1
X_4015_ clknet_leaf_19_wb_clk_i _0503_ net285 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2492__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout134_X net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4655__424 vssd1 vssd1 vccd1 vccd1 _4655__424/HI net424 sky130_fd_sc_hd__conb_1
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4192__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2483__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_44_Left_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2214__B net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2130_ net214 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0930_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_53_Left_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2061_ team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] net112 net138 net663 vssd1
+ vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3423__C1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2963_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] net163 _1483_ net216
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[10\]
+ sky130_fd_sc_hd__o22a_1
X_1914_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] vssd1 vssd1 vccd1 vccd1
+ _0837_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_62_Left_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2894_ net157 net151 vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__nand2_1
X_4639__408 vssd1 vssd1 vccd1 vccd1 _4639__408/HI net408 sky130_fd_sc_hd__conb_1
X_4633_ net402 vssd1 vssd1 vccd1 vccd1 la_data_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_53_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4564_ net440 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3515_ net246 vssd1 vssd1 vccd1 vccd1 _0047_ sky130_fd_sc_hd__inv_2
XANTENNA__4065__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4495_ net307 vssd1 vssd1 vccd1 vccd1 ADR_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3446_ team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] _1715_ _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[13\]
+ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__a22o_1
X_3377_ team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] net180 net179 team_10_WB.instance_to_wrap.dispFSM.guesses\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2328_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[5\] _0858_ vssd1 vssd1
+ vccd1 vccd1 _1104_ sky130_fd_sc_hd__xor2_1
X_2259_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0798_ _1036_ _1037_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_28_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1976__C1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4408__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1991__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2940__A1 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input24_A wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4088__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3300_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] _0817_ vssd1 vssd1 vccd1
+ vccd1 _1681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4280_ clknet_leaf_16_wb_clk_i _0670_ _0269_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3231_ _1637_ _1611_ _1636_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__and3b_1
X_3162_ _0812_ net4 _0906_ _1582_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__and4_1
XFILLER_0_55_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2113_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__nand2b_1
X_3093_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net198 vssd1 vssd1 vccd1
+ vccd1 _1541_ sky130_fd_sc_hd__and2_1
X_2044_ team_10_WB.instance_to_wrap.dispFSM.guesses\[68\] net115 net136 net674 vssd1
+ vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3995_ clknet_leaf_24_wb_clk_i _0485_ _0063_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3411__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2946_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[0\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[2\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[3\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\]
+ net165 vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__a41o_1
XANTENNA__2135__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2877_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[2\] _1461_ vssd1 vssd1 vccd1
+ vccd1 _1462_ sky130_fd_sc_hd__mux2_1
X_4616_ net388 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XFILLER_0_44_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1973__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4547_ net359 vssd1 vssd1 vccd1 vccd1 DAT_O[21] sky130_fd_sc_hd__buf_2
X_4478_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[35\]
+ _0461_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3429_ net303 team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _0815_ net211 vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_55_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout299_X net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3478__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2438__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2989__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4380__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1964__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3948__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3469__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2429__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2800_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\] team_10_WB.instance_to_wrap.lcdPlayer.currentState\[4\]
+ _1403_ vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__mux2_1
X_3780_ net291 vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2731_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ _1356_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4401_ clknet_leaf_6_wb_clk_i _0786_ _0384_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2662_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ _1318_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2593_ _0910_ _1276_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4332_ clknet_leaf_19_wb_clk_i net628 _0321_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\]
+ sky130_fd_sc_hd__dfrtp_1
X_4571__447 vssd1 vssd1 vccd1 vccd1 net447 _4571__447/LO sky130_fd_sc_hd__conb_1
X_4263_ clknet_leaf_4_wb_clk_i _0653_ _0252_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.correct\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout219 team_10_WB.instance_to_wrap.gamelogic.state\[0\] vssd1 vssd1 vccd1 vccd1
+ net219 sky130_fd_sc_hd__buf_2
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
X_3214_ _1626_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4103__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4194_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[56\]
+ _0183_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[56\] sky130_fd_sc_hd__dfrtp_1
X_3145_ _1569_ _1573_ _1574_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__and3_1
X_3076_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] _1532_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[74\] sky130_fd_sc_hd__mux2_1
X_2027_ _0888_ _0908_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3978_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[15\]
+ _0046_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2929_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] net151 net120 net647
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[34\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_57_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold262 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\] vssd1 vssd1 vccd1
+ vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\] vssd1 vssd1 vccd1
+ vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\] vssd1 vssd1 vccd1
+ vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 net82 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3084__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1879__A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2898__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4126__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4276__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 wbs_adr_i[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__buf_1
Xclkbuf_2_0__f_wb_clk_i clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_2_0__leaf_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3340__Y _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3901_ net247 vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3090__A3 net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3832_ net257 vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3763_ net271 vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__inv_2
X_2714_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ _1347_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__and3_1
X_3694_ net233 vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__inv_2
X_2645_ net1 net157 team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 _1307_ sky130_fd_sc_hd__and3b_1
XFILLER_0_61_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4401__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4315_ clknet_leaf_20_wb_clk_i _0705_ _0304_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[38\]
+ sky130_fd_sc_hd__dfstp_1
X_2576_ net221 net227 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] vssd1
+ vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4246_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[2\]
+ _0235_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4177_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[2\]
+ _0166_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2105__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128_ _1286_ _1288_ _1291_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__or4b_1
X_3059_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__B2 team_10_WB.instance_to_wrap.host_row2\[74\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4149__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_670 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3057__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_776 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4221__Q team_10_WB.instance_to_wrap.host_row2\[83\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2430_ _0993_ _1185_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__and2_2
XANTENNA__3335__Y _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_11 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2361_ _1096_ _1131_ _1135_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__and3_1
X_4100_ clknet_leaf_12_wb_clk_i _0571_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2292_ _0842_ _0866_ _1070_ _0865_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__o22a_1
X_4031_ clknet_leaf_11_wb_clk_i _0516_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3815_ net255 vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
X_3746_ net295 vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4441__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3677_ net240 vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__inv_2
XANTENNA__2430__X _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2797__B net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2628_ _0009_ _0010_ _0008_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[0\]
+ sky130_fd_sc_hd__or3_1
X_2559_ net219 _0952_ _1024_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4229_ clknet_leaf_0_wb_clk_i _0645_ _0218_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2798__C1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_795 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2014__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4314__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1930_ net226 _0851_ vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4464__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput11 wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_2
X_3600_ net262 vssd1 vssd1 vccd1 vccd1 _0132_ sky130_fd_sc_hd__inv_2
X_4580_ net201 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput22 wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 wbs_adr_i[3] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3531_ net269 vssd1 vssd1 vccd1 vccd1 _0063_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3462_ team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] net171 _1833_ _1835_ vssd1
+ vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3393_ team_10_WB.instance_to_wrap.host_row2\[83\] net173 net167 team_10_WB.instance_to_wrap.host_row2\[75\]
+ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__a221o_1
X_2413_ _1167_ _1173_ _1174_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2344_ _0823_ _1857_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] vssd1 vssd1
+ vccd1 vccd1 _1120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4533__345 vssd1 vssd1 vccd1 vccd1 _4533__345/HI net345 sky130_fd_sc_hd__conb_1
X_2275_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] _1056_ vssd1 vssd1
+ vccd1 vccd1 _1057_ sky130_fd_sc_hd__nor2_1
X_4014_ clknet_leaf_25_wb_clk_i _0502_ net273 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_36_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_954 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3729_ net236 vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2235__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1994__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_724 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4517__329 vssd1 vssd1 vccd1 vccd1 _4517__329/HI net329 sky130_fd_sc_hd__conb_1
X_2060_ team_10_WB.instance_to_wrap.dispFSM.guesses\[52\] net109 net135 net633 vssd1
+ vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_707 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2962_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\] net161 _1483_ net217 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[9\] sky130_fd_sc_hd__o22a_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1913_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\] vssd1 vssd1 vccd1 vccd1
+ _0836_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4632_ net401 vssd1 vssd1 vccd1 vccd1 la_data_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2893_ net166 net156 vssd1 vssd1 vccd1 vccd1 _1472_ sky130_fd_sc_hd__nor2_1
X_4604__379 vssd1 vssd1 vccd1 vccd1 _4604__379/HI net379 sky130_fd_sc_hd__conb_1
XFILLER_0_53_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4563_ net375 vssd1 vssd1 vccd1 vccd1 WE_O sky130_fd_sc_hd__buf_2
X_4494_ net306 vssd1 vssd1 vccd1 vccd1 ADR_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3514_ net246 vssd1 vssd1 vccd1 vccd1 _0046_ sky130_fd_sc_hd__inv_2
X_3445_ net232 _1819_ _1817_ _1812_ _1807_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3376_ team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] net174 net171 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\]
+ _1753_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2327_ team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\] _0854_ vssd1 vssd1
+ vccd1 vccd1 _1103_ sky130_fd_sc_hd__xnor2_1
X_2258_ team_10_WB.instance_to_wrap.gamelogic.setWord\[39\] _0798_ _0799_ team_10_WB.instance_to_wrap.gamelogic.setWord\[38\]
+ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout289_A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2189_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] net213 vssd1 vssd1 vccd1
+ vccd1 _0978_ sky130_fd_sc_hd__nand2_1
XANTENNA__3398__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3414__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_X net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2940__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input17_A wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2456__B2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3405__B1 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2241__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2392__A0 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3230_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ _1633_ vssd1 vssd1 vccd1 vccd1 _1637_ sky130_fd_sc_hd__and3_1
X_3161_ team_10_WB.instance_to_wrap.dispFSM.msg\[2\] _0886_ _1274_ _1581_ _1589_ vssd1
+ vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__o32a_1
X_2112_ team_10_WB.instance_to_wrap.dispFSM.guesses\[0\] net114 net141 net704 vssd1
+ vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3092_ net204 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] net187 _1540_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[82\] sky130_fd_sc_hd__a31o_1
X_2043_ team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] net143 net107 net582 vssd1
+ vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_941 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4032__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3994_ clknet_leaf_24_wb_clk_i _0484_ _0062_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_col\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] net126 _1474_ vssd1
+ vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2876_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] net224 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__or3b_1
X_4498__310 vssd1 vssd1 vccd1 vccd1 _4498__310/HI net310 sky130_fd_sc_hd__conb_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4615_ team_10_WB.instance_to_wrap.gamelogic.red vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_1
XANTENNA__2422__Y _1184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4546_ net358 vssd1 vssd1 vccd1 vccd1 DAT_O[20] sky130_fd_sc_hd__buf_2
XANTENNA__4182__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2151__A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4539__351 vssd1 vssd1 vccd1 vccd1 _4539__351/HI net351 sky130_fd_sc_hd__conb_1
XANTENNA_fanout204_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4477_ clknet_leaf_4_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[34\]
+ _0460_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
X_3428_ team_10_WB.instance_to_wrap.host_row1\[53\] net302 _1699_ vssd1 vssd1 vccd1
+ vccd1 _1803_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ team_10_WB.instance_to_wrap.host_row1\[41\] _1693_ _1703_ team_10_WB.instance_to_wrap.host_row1\[65\]
+ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__a221o_1
XANTENNA__3332__C1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_X net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2211__D net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3444__X _1819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2126__A0 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3620__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4055__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_454 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2730_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ team_10_WB.instance_to_wrap.clock_div.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__a21oi_1
X_2661_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\] _1319_ vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[0\] sky130_fd_sc_hd__and2b_1
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4400_ clknet_leaf_1_wb_clk_i _0785_ _0383_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2592_ _0910_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__and2_1
X_4331_ clknet_leaf_20_wb_clk_i _0721_ _0320_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[54\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4262_ clknet_leaf_1_wb_clk_i _0652_ _0251_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout209 team_10_WB.instance_to_wrap.hostdisp.Cstate vssd1 vssd1 vccd1 vccd1 net209
+ sky130_fd_sc_hd__buf_2
X_3213_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\] _1621_ vssd1 vssd1 vccd1 vccd1
+ _1626_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4193_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[55\]
+ _0182_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[55\] sky130_fd_sc_hd__dfrtp_1
X_3144_ _1557_ _1571_ _1572_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3075_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__mux2_1
XANTENNA__3530__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2026_ _0888_ _0908_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout154_A net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3977_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[14\]
+ _0045_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1985__A team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2928_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] net154 net123 net651
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[33\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3396__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2859_ _1450_ _1451_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[6\]
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_57_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4529_ net341 vssd1 vssd1 vccd1 vccd1 DAT_O[3] sky130_fd_sc_hd__buf_2
Xhold230 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\] vssd1 vssd1 vccd1
+ vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold241 team_10_WB.instance_to_wrap.dispFSM.guesses\[44\] vssd1 vssd1 vccd1 vccd1
+ net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[26\] vssd1 vssd1 vccd1
+ vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 team_10_WB.instance_to_wrap.host_row1\[75\] vssd1 vssd1 vccd1 vccd1 net720
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3705__A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 team_10_WB.instance_to_wrap.clock_div.count\[8\] vssd1 vssd1 vccd1 vccd1
+ net731 sky130_fd_sc_hd__dlygate4sd3_1
X_4617__389 vssd1 vssd1 vccd1 vccd1 _4617__389/HI net389 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_5_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3320__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3387__A2 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_800 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_833 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput9 wbs_adr_i[10] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_1
XFILLER_0_8_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ net264 vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3831_ net260 vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3762_ net295 vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__inv_2
XANTENNA__3378__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2713_ net556 _1347_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[4\]
+ sky130_fd_sc_hd__xor2_1
X_3693_ net233 vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__inv_2
X_2644_ _0923_ _0947_ _1302_ _0924_ _0922_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[3\]
+ sky130_fd_sc_hd__a32o_1
X_2575_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[2\] net227 net221 vssd1
+ vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2889__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4314_ clknet_leaf_25_wb_clk_i _0704_ _0303_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4220__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4245_ clknet_leaf_30_wb_clk_i net534 _0234_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4176_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[1\]
+ _0165_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__dfrtp_1
X_3127_ _1862_ _1555_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] vssd1
+ vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__a21o_1
XANTENNA__4370__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3058_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _1523_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\] sky130_fd_sc_hd__mux2_1
XANTENNA__2147__Y _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2009_ team_10_WB.instance_to_wrap.keypadplayer.scan_col\[3\] team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\]
+ net222 net223 vssd1 vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__nor4_2
XANTENNA_fanout157_X net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_744 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2360_ _1124_ _1134_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_23 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2291_ net5 _0844_ net196 vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__and3_1
XANTENNA__4393__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ clknet_leaf_10_wb_clk_i _0515_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_25 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2559__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2424__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ net247 vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_755 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3745_ net280 vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3676_ net277 vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout117_A net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2627_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\] _1074_ _1297_ vssd1 vssd1
+ vccd1 vccd1 _0008_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_7_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2558_ _1243_ _1247_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__nor2_1
X_2489_ net499 net129 _1189_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1
+ vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4228_ clknet_leaf_0_wb_clk_i _0644_ _0217_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout274_X net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4159_ clknet_leaf_28_wb_clk_i _0628_ _0148_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4116__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2486__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 wbs_adr_i[13] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
Xinput34 wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput23 wbs_adr_i[23] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
X_3530_ net269 vssd1 vssd1 vccd1 vccd1 _0062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3461_ team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] net181 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__a221o_1
X_3392_ team_10_WB.instance_to_wrap.host_row1\[75\] _1708_ net180 team_10_WB.instance_to_wrap.host_row2\[59\]
+ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__a22o_1
X_2412_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[9\]
+ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2343_ _0870_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2274_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0800_ _1051_ _1052_ _1049_
+ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4013_ clknet_leaf_19_wb_clk_i _0501_ net273 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4139__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2419__A net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2492__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4289__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3441__B2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3441__A1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout234_A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__A1_N team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3944__RESET_B _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1989_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] net147 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[10\]
+ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2952__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3728_ net234 vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__inv_2
X_3659_ net282 vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3713__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2483__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2235__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1994__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1994__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_736 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4556__368 vssd1 vssd1 vccd1 vccd1 _4556__368/HI net368 sky130_fd_sc_hd__conb_1
XANTENNA__3623__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2459__C1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4431__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4227__Q team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2474__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3423__A1 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_655 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2961_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] net163 _1483_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[8\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1912_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[23\] vssd1 vssd1 vccd1 vccd1
+ _0835_ sky130_fd_sc_hd__inv_2
X_4631_ net400 vssd1 vssd1 vccd1 vccd1 la_data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_57_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2892_ net193 _1471_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[7\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4500__312 vssd1 vssd1 vccd1 vccd1 _4500__312/HI net312 sky130_fd_sc_hd__conb_1
X_4562_ net374 vssd1 vssd1 vccd1 vccd1 STB_O sky130_fd_sc_hd__buf_2
XFILLER_0_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4493_ net305 vssd1 vssd1 vccd1 vccd1 ADR_O[0] sky130_fd_sc_hd__buf_2
X_3513_ net246 vssd1 vssd1 vccd1 vccd1 _0045_ sky130_fd_sc_hd__inv_2
XANTENNA__2934__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3444_ team_10_WB.instance_to_wrap.host_row2\[45\] net174 net169 team_10_WB.instance_to_wrap.host_row1\[61\]
+ _1818_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3375_ team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] net168 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__a22o_1
XANTENNA__2162__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload19_A clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2326_ _1100_ _1101_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nand2_1
X_2257_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net217 vssd1 vssd1 vccd1
+ vccd1 _1039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2188_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net216 vssd1 vssd1 vccd1
+ vccd1 _0977_ sky130_fd_sc_hd__nand2_1
X_4661__430 vssd1 vssd1 vccd1 vccd1 _4661__430/HI net430 sky130_fd_sc_hd__conb_1
XANTENNA__3414__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2925__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4454__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__B net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2456__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Left_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2208__A2 _0995_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_647 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3341__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3160_ _0903_ _1588_ net195 vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__o21a_1
X_3091_ team_10_WB.instance_to_wrap.gamelogic.setWord\[34\] net198 vssd1 vssd1 vccd1
+ vccd1 _1540_ sky130_fd_sc_hd__and2_1
X_2111_ team_10_WB.instance_to_wrap.dispFSM.guesses\[1\] net110 net137 net660 vssd1
+ vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__o22a_1
Xhold1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe vssd1 vssd1 vccd1 vccd1
+ net458 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2042_ team_10_WB.instance_to_wrap.dispFSM.guesses\[70\] net111 net138 net672 vssd1
+ vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4645__414 vssd1 vssd1 vccd1 vccd1 _4645__414/HI net414 sky130_fd_sc_hd__conb_1
XFILLER_0_58_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2416__B net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3971__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3993_ clknet_leaf_25_wb_clk_i _0483_ _0061_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe
+ sky130_fd_sc_hd__dfrtp_1
X_2944_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[4\] _0831_ net165 vssd1 vssd1
+ vccd1 vccd1 _1475_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2875_ net193 _1460_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[1\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__2432__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4614_ team_10_WB.instance_to_wrap.gamelogic.green vssd1 vssd1 vccd1 vccd1 net73
+ sky130_fd_sc_hd__clkbuf_1
X_4545_ net357 vssd1 vssd1 vccd1 vccd1 DAT_O[19] sky130_fd_sc_hd__buf_2
XANTENNA__2907__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4476_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[33\]
+ _0459_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3427_ team_10_WB.instance_to_wrap.host_row2\[61\] team_10_WB.instance_to_wrap.dispFSM.guesses\[37\]
+ net301 vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_X clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ team_10_WB.instance_to_wrap.host_row2\[41\] net174 net173 team_10_WB.instance_to_wrap.host_row2\[81\]
+ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_0_wb_clk_i_X clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2309_ net693 _1076_ _1077_ net160 vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__a31o_1
X_3289_ _1672_ _1673_ vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2438__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3020__C1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_374 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2429__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3994__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2660_ _1307_ _1310_ _1313_ _1317_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_41_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2591_ _0908_ _1219_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4330_ clknet_leaf_19_wb_clk_i _0720_ _0319_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_4261_ clknet_leaf_4_wb_clk_i _0651_ _0250_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.red
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3212_ net726 _1622_ _1625_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4192_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[54\]
+ _0181_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[54\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3143_ _1557_ _1572_ _1571_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__o21ai_1
X_3074_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] _1531_ net207 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[73\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2427__A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2025_ net3 _0901_ _0907_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_59_Left_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3976_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[13\]
+ _0044_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout147_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2927_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] net152 net120 net659
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[32\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__2053__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2858_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\] _1448_ net176
+ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__o21ai_1
XANTENNA__4150__Q net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2789_ _1393_ _1395_ _1396_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__nor4_1
Xhold220 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[42\] vssd1 vssd1 vccd1
+ vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ net340 vssd1 vssd1 vccd1 vccd1 DAT_O[2] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] vssd1 vssd1 vccd1 vccd1
+ net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 team_10_WB.instance_to_wrap.dispFSM.guesses\[26\] vssd1 vssd1 vccd1 vccd1
+ net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] vssd1 vssd1 vccd1 vccd1
+ net710 sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[16\]
+ _0442_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
Xhold264 team_10_WB.instance_to_wrap.dispFSM.guesses\[10\] vssd1 vssd1 vccd1 vccd1
+ net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold275 team_10_WB.instance_to_wrap.clock_div.count\[20\] vssd1 vssd1 vccd1 vccd1
+ net732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3721__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2898__A2 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_845 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4172__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3830_ net259 vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3761_ net292 vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2712_ _1347_ _1348_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[3\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3692_ net284 vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__inv_2
X_2643_ _0953_ _1306_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[2\]
+ sky130_fd_sc_hd__or2_1
X_2574_ net222 net227 vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4313_ clknet_leaf_12_wb_clk_i _0703_ _0302_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3017__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4244_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[0\]
+ _0233_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4175_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[0\]
+ _0164_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__dfrtp_1
X_3126_ _1286_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__nor3_1
XANTENNA__2428__Y _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3057_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout264_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2008_ net222 _0890_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3959_ clknet_leaf_27_wb_clk_i _0010_ _0027_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4045__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4195__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_35 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2290_ _0842_ _1067_ _0859_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ net273 vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_26 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2424__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ net298 vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3675_ net242 vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_31_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2626_ _0828_ _1117_ _1132_ _1235_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3536__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2557_ _1239_ _1241_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__a21oi_1
X_2488_ net518 net130 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[6\] vssd1
+ vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4227_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.host_message_reg.next_state
+ _0216_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.Cstate
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_39_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4158_ clknet_leaf_28_wb_clk_i net459 _0147_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge
+ sky130_fd_sc_hd__dfrtp_1
X_4089_ clknet_leaf_13_wb_clk_i _0560_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3109_ team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked _0893_ net227 vssd1 vssd1
+ vccd1 vccd1 _1548_ sky130_fd_sc_hd__and3_2
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2014__A3 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2486__B1 net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2238__B1 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_859 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4210__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
Xinput35 wbs_adr_i[5] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 wbs_adr_i[24] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4360__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2260__A team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2961__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3460_ team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] net175 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[78\]
+ _0821_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__a221o_1
X_3391_ team_10_WB.instance_to_wrap.host_row2\[51\] net170 _1703_ team_10_WB.instance_to_wrap.host_row1\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__a22o_1
X_2411_ team_10_WB.instance_to_wrap.clock_div.count\[11\] team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__or4b_1
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2342_ _0820_ _0864_ _0842_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2273_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _0798_ _0801_ team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__o22a_1
X_4012_ clknet_leaf_19_wb_clk_i _0500_ net285 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2477__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2419__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3030__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2435__A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__o22a_1
X_3727_ net234 vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__inv_2
XANTENNA__2952__B2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3658_ net247 vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2609_ _0886_ _1274_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nor2_2
X_3589_ net268 vssd1 vssd1 vccd1 vccd1 _0121_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3432__A2 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4383__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3463__X _1837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout190 net192 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2459__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4567__443 vssd1 vssd1 vccd1 vccd1 net443 _4567__443/LO sky130_fd_sc_hd__conb_1
XANTENNA_clkload5_A clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3423__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ net126 _1482_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__nand2_2
XFILLER_0_57_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2891_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] net1 _1227_ vssd1 vssd1 vccd1
+ vccd1 _1471_ sky130_fd_sc_hd__mux2_1
X_1911_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\] vssd1 vssd1 vccd1 vccd1
+ _0834_ sky130_fd_sc_hd__inv_2
X_4630_ net399 vssd1 vssd1 vccd1 vccd1 la_data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_56_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4561_ net373 vssd1 vssd1 vccd1 vccd1 SEL_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_350 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4492_ clknet_leaf_14_wb_clk_i _0017_ _0475_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfrtp_1
X_3512_ net250 vssd1 vssd1 vccd1 vccd1 _0044_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_wb_clk_i_X clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3443_ team_10_WB.instance_to_wrap.host_row2\[53\] net170 net167 team_10_WB.instance_to_wrap.host_row2\[77\]
+ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__a22o_1
XANTENNA__4106__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3374_ _1747_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__or3_2
XANTENNA__3025__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2325_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\]
+ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1858_ vssd1 vssd1 vccd1 vccd1
+ _1101_ sky130_fd_sc_hd__or4b_1
X_2256_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net217 vssd1 vssd1 vccd1
+ vccd1 _1038_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_25_Left_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout177_A net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2187_ team_10_WB.instance_to_wrap.gamelogic.setWord\[10\] net216 vssd1 vssd1 vccd1
+ vccd1 _0976_ sky130_fd_sc_hd__or2_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3414__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_731 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1976__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3724__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3102__A1 net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4523__335 vssd1 vssd1 vccd1 vccd1 _4523__335/HI net335 sky130_fd_sc_hd__conb_1
XFILLER_0_54_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3169__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4129__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1922__A_N net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4279__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3090_ net207 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[41\] net190 _1539_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[81\] sky130_fd_sc_hd__a31o_1
X_2110_ team_10_WB.instance_to_wrap.dispFSM.guesses\[2\] net112 net141 net721 vssd1
+ vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__o22a_1
Xhold2 team_10_WB.instance_to_wrap.keypadFSMHost.strobe vssd1 vssd1 vccd1 vccd1 net459
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2041_ net595 net144 net108 net611 vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__a22o_1
X_4610__385 vssd1 vssd1 vccd1 vccd1 _4610__385/HI net385 sky130_fd_sc_hd__conb_1
X_3992_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[29\]
+ _0060_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2943_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] net158 vssd1 vssd1 vccd1
+ vccd1 _1474_ sky130_fd_sc_hd__nand2_1
X_2874_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[1\] _1459_ vssd1 vssd1 vccd1
+ vccd1 _1460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4613_ team_10_WB.instance_to_wrap.blue vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_1
X_4544_ net356 vssd1 vssd1 vccd1 vccd1 DAT_O[18] sky130_fd_sc_hd__buf_2
XFILLER_0_40_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[32\]
+ _0458_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3426_ team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.dispFSM.guesses\[69\]
+ net302 vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3357_ team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] net170 net169 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ _1735_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__a221o_1
X_2308_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] _1078_ _1083_
+ _1082_ _1079_ vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__o32a_1
X_3288_ net635 _1671_ net231 vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__o21ai_1
X_2239_ _0796_ net212 _0799_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _1020_
+ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4507__319 vssd1 vssd1 vccd1 vccd1 _4507__319/HI net319 sky130_fd_sc_hd__conb_1
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4421__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input22_A wbs_adr_i[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_924 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_158 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_180 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2590_ net195 _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4260_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[3\]
+ _0249_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_3211_ net172 _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__nor2_1
X_4191_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[53\]
+ _0180_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[53\] sky130_fd_sc_hd__dfrtp_1
X_3142_ _1286_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__and3b_1
XFILLER_0_24_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3073_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\]
+ net191 vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2024_ _0904_ _0906_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3975_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[12\]
+ _0043_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3539__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3098__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2926_ net613 net156 net125 net643 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[31\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__4444__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2857_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[6\] _1448_ vssd1 vssd1
+ vccd1 vccd1 _1450_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2788_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1397_ vssd1 vssd1 vccd1 vccd1
+ _1398_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold210 team_10_WB.instance_to_wrap.clock_div.count\[3\] vssd1 vssd1 vccd1 vccd1
+ net667 sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ net339 vssd1 vssd1 vccd1 vccd1 DAT_O[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold243 team_10_WB.instance_to_wrap.dispFSM.guesses\[25\] vssd1 vssd1 vccd1 vccd1
+ net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold232 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1
+ net689 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 team_10_WB.instance_to_wrap.dispFSM.guesses\[77\] vssd1 vssd1 vccd1 vccd1
+ net678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\] vssd1 vssd1 vccd1
+ vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\] vssd1 vssd1 vccd1 vccd1
+ net733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] vssd1 vssd1 vccd1 vccd1
+ net711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[15\]
+ _0441_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3409_ team_10_WB.instance_to_wrap.host_row1\[44\] _1693_ net173 team_10_WB.instance_to_wrap.host_row2\[84\]
+ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__a22o_1
X_4389_ clknet_leaf_3_wb_clk_i _0774_ _0372_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_5_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3961__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4317__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2528__A _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4529__341 vssd1 vssd1 vccd1 vccd1 _4529__341/HI net341 sky130_fd_sc_hd__conb_1
XANTENNA__4467__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3760_ net293 vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2711_ net667 _1345_ vssd1 vssd1 vccd1 vccd1 _1348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3691_ net284 vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2642_ net219 _0952_ _1306_ _0951_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2573_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[3\] _1257_ vssd1 vssd1
+ vccd1 vccd1 _1258_ sky130_fd_sc_hd__xnor2_1
X_4312_ clknet_leaf_16_wb_clk_i _0702_ _0301_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4243_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[7\]
+ _0232_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4174_ clknet_leaf_26_wb_clk_i _0643_ _0163_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3125_ _0824_ _1861_ _1555_ _1291_ vssd1 vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a31o_1
XANTENNA__3033__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3056_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] _1522_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\] sky130_fd_sc_hd__mux2_2
X_2007_ net220 net221 vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__or2_1
XANTENNA__2274__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3471__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3958_ clknet_leaf_27_wb_clk_i _0009_ _0026_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_2909_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\] net155 net122 net680
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[14\]
+ sky130_fd_sc_hd__o22a_1
X_3889_ net279 vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_X net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4630__399 vssd1 vssd1 vccd1 vccd1 _4630__399/HI net399 sky130_fd_sc_hd__conb_1
XFILLER_0_49_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3453__B1 net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3089__A team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3812_ net287 vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__inv_2
XANTENNA_27 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3743_ net280 vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3674_ net248 vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__inv_2
Xoutput101 net184 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2625_ _0010_ _0007_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[1\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2556_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] _1243_ _1245_
+ _1242_ _1239_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__o221a_1
X_2487_ net525 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1
+ vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__a22o_1
X_4226_ clknet_leaf_11_wb_clk_i net439 _0215_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4157_ clknet_leaf_28_wb_clk_i net461 _0146_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge1
+ sky130_fd_sc_hd__dfrtp_1
X_3108_ net730 net40 net42 vssd1 vssd1 vccd1 vccd1 _0017_ sky130_fd_sc_hd__and3b_1
X_4088_ clknet_leaf_12_wb_clk_i _0559_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3039_ team_10_WB.instance_to_wrap.gamelogic.setWord\[16\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1514_ sky130_fd_sc_hd__mux2_1
XANTENNA__3444__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2798__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2014__A4 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4012__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4162__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2806__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2238__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1997__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput36 wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_1
Xinput14 wbs_adr_i[15] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2260__B _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2410_ team_10_WB.instance_to_wrap.clock_div.count\[2\] team_10_WB.instance_to_wrap.clock_div.count\[4\]
+ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__or3_1
X_3390_ _1763_ _1765_ _1766_ net303 vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__o31a_1
X_2341_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\] _1112_ _1115_ vssd1 vssd1
+ vccd1 vccd1 _1117_ sky130_fd_sc_hd__and3b_1
X_2272_ _0792_ net215 _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] vssd1
+ vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__a22o_1
XANTENNA__3091__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4011_ clknet_leaf_19_wb_clk_i _0499_ net285 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[3\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_36_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3426__A0 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4035__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1988__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2435__B _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1987_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net150 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout122_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3547__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4185__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3726_ net234 vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__inv_2
X_3657_ net263 vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2165__A0 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\] _1275_ _1284_ _1289_
+ vssd1 vssd1 vccd1 vccd1 _0014_ sky130_fd_sc_hd__a22o_1
X_3588_ net267 vssd1 vssd1 vccd1 vccd1 _0120_ sky130_fd_sc_hd__inv_2
X_2539_ team_10_WB.instance_to_wrap.host_col\[3\] _0852_ _1179_ vssd1 vssd1 vccd1
+ vccd1 _0487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4209_ clknet_leaf_18_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\]
+ _0198_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[71\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1979__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_2
Xfanout180 _1709_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_4
XANTENNA__2459__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4058__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3408__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2255__B net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1910_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\] vssd1 vssd1 vccd1 vccd1
+ _0833_ sky130_fd_sc_hd__inv_2
X_2890_ net193 _1470_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[6\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4560_ net372 vssd1 vssd1 vccd1 vccd1 SEL_O[2] sky130_fd_sc_hd__buf_2
XFILLER_0_53_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3511_ net250 vssd1 vssd1 vccd1 vccd1 _0043_ sky130_fd_sc_hd__inv_2
XANTENNA__2934__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4491_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_state _0474_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.Cstate sky130_fd_sc_hd__dfrtp_1
X_3442_ _1800_ _1813_ _1815_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3373_ team_10_WB.instance_to_wrap.host_row1\[66\] _1703_ net180 team_10_WB.instance_to_wrap.host_row2\[58\]
+ _1748_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__a221o_1
X_2324_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__nor2_1
X_2255_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net215 vssd1 vssd1 vccd1
+ vccd1 _1037_ sky130_fd_sc_hd__or2_1
X_2186_ _0822_ _0952_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_62_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_668 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout125_X net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4689_ net183 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_1
X_3709_ net235 vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2138__A0 team_10_WB.instance_to_wrap.gamelogic.letter\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4200__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4350__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4562__374 vssd1 vssd1 vccd1 vccd1 _4562__374/HI net374 sky130_fd_sc_hd__conb_1
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2916__A2 _1181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3326__C1 _1705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3341__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold3 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge vssd1 vssd1 vccd1 vccd1
+ net460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2040_ team_10_WB.instance_to_wrap.dispFSM.guesses\[72\] net113 net140 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__o22a_1
XANTENNA__2266__A team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3991_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[28\]
+ _0059_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2942_ net212 net156 net125 net602 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[47\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net224 vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__or3b_1
XANTENNA__3097__A team_10_WB.instance_to_wrap.gamelogic.setWord\[37\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4612_ net387 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
X_4543_ net355 vssd1 vssd1 vccd1 vccd1 DAT_O[17] sky130_fd_sc_hd__buf_2
XANTENNA__2907__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4474_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[31\]
+ _0457_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4223__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload24_A clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3036__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3425_ team_10_WB.instance_to_wrap.host_row1\[45\] net302 _1693_ vssd1 vssd1 vccd1
+ vccd1 _1800_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2032__B1_N net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3332__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3356_ team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] net167 _1732_ _1734_ vssd1
+ vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__a211o_1
X_3287_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[17\] _1671_ vssd1 vssd1 vccd1
+ vccd1 _1672_ sky130_fd_sc_hd__and2_1
X_2307_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2238_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _0804_ _0800_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4373__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3096__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2169_ team_10_WB.instance_to_wrap.correct\[0\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4546__358 vssd1 vssd1 vccd1 vccd1 _4546__358/HI net358 sky130_fd_sc_hd__conb_1
XFILLER_0_49_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input15_A wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4396__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4651__420 vssd1 vssd1 vccd1 vccd1 _4651__420/HI net420 sky130_fd_sc_hd__conb_1
X_4190_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[52\]
+ _0179_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[52\] sky130_fd_sc_hd__dfrtp_1
X_3210_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ _1621_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3141_ _1563_ _1570_ _0905_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] _1530_ net204 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[72\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2023_ _0893_ _0895_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_18_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3974_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[11\]
+ _0042_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_2925_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\] net154 net122 net648
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[30\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2443__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2856_ _1448_ _1449_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[5\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2787_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__and4b_1
XANTENNA__3002__B2 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold211 team_10_WB.instance_to_wrap.dispFSM.guesses\[50\] vssd1 vssd1 vccd1 vccd1
+ net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 team_10_WB.instance_to_wrap.dispFSM.guesses\[66\] vssd1 vssd1 vccd1 vccd1
+ net657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3555__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4526_ net338 vssd1 vssd1 vccd1 vccd1 DAT_O[0] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_57_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold244 team_10_WB.instance_to_wrap.dispFSM.guesses\[28\] vssd1 vssd1 vccd1 vccd1
+ net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 team_10_WB.instance_to_wrap.host_row1\[48\] vssd1 vssd1 vccd1 vccd1 net679
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A net209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold233 team_10_WB.instance_to_wrap.dispFSM.guesses\[30\] vssd1 vssd1 vccd1 vccd1
+ net690 sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[14\]
+ _0440_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xhold277 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\] vssd1 vssd1 vccd1
+ vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\] vssd1 vssd1 vccd1 vccd1
+ net723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold255 team_10_WB.instance_to_wrap.dispFSM.guesses\[73\] vssd1 vssd1 vccd1 vccd1
+ net712 sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ team_10_WB.instance_to_wrap.host_row1\[52\] _1699_ net167 team_10_WB.instance_to_wrap.host_row2\[76\]
+ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4388_ clknet_leaf_6_wb_clk_i _0773_ _0371_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_input7_A wb_rst_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3339_ _1687_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4119__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2044__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635__404 vssd1 vssd1 vccd1 vccd1 _4635__404/HI net404 sky130_fd_sc_hd__conb_1
XFILLER_0_47_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2809__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4681__435 vssd1 vssd1 vccd1 vccd1 _4681__435/HI net435 sky130_fd_sc_hd__conb_1
XFILLER_0_54_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_700 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4181__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2710_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ net235 vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__inv_2
X_2641_ _0945_ _1305_ _0936_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__a21o_1
X_2572_ net220 net227 vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4311_ clknet_leaf_16_wb_clk_i _0701_ _0300_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4242_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[6\]
+ _0231_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4173_ clknet_leaf_25_wb_clk_i _0642_ _0162_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_2_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3124_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__nor2_1
X_3055_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[24\]
+ net187 vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__mux2_1
XANTENNA__2259__C1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2006_ net220 team_10_WB.instance_to_wrap.keypadplayer.scan_col\[2\] vssd1 vssd1
+ vccd1 vccd1 _0889_ sky130_fd_sc_hd__nor2_1
XANTENNA__4411__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2274__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3957_ clknet_leaf_27_wb_clk_i _0008_ _0025_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2908_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[21\] _1181_ _1472_ net616
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3888_ net275 vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2839_ _0518_ _1439_ _1436_ _1411_ vssd1 vssd1 vccd1 vccd1 _0003_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4509_ net321 vssd1 vssd1 vccd1 vccd1 ADR_O[16] sky130_fd_sc_hd__buf_2
XANTENNA__2635__Y _1302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_9_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4434__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_346 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3089__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ net273 vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
XANTENNA_28 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4262__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3742_ net293 vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3673_ net263 vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2624_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\] _1074_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0007_ sky130_fd_sc_hd__a22o_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[3] sky130_fd_sc_hd__buf_2
XANTENNA__2192__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2555_ _1246_ _1239_ _1244_ vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__and3b_1
X_2486_ net679 net130 net126 team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] _1190_
+ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4225_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[87\]
+ _0214_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[87\] sky130_fd_sc_hd__dfrtp_1
X_4156_ clknet_leaf_23_wb_clk_i _0627_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked
+ sky130_fd_sc_hd__dfrtp_1
X_3107_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1395_ _1547_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.lcd_en sky130_fd_sc_hd__nor3_1
XFILLER_0_37_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4087_ clknet_leaf_12_wb_clk_i _0558_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4664__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2247__A2 net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3038_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] _1513_ net208 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[55\] sky130_fd_sc_hd__mux2_1
XANTENNA_fanout155_X net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2184__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2955__B1 net159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4457__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2486__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1997__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2822__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 wbs_adr_i[7] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 wbs_adr_i[16] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
Xinput26 wbs_adr_i[26] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3371__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2340_ _1112_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__nand2_1
XANTENNA__2269__A team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2271_ team_10_WB.instance_to_wrap.gamelogic.setWord\[26\] _0803_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ _1048_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__o221a_1
X_4010_ clknet_leaf_25_wb_clk_i _0498_ net273 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__2477__A2 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2229__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] _0874_ _0882_ net159 vssd1
+ vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_60_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2937__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3725_ net244 vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3656_ net271 vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__inv_2
X_2607_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\] team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\]
+ _1288_ _1270_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__or4b_1
XFILLER_0_11_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3587_ net253 vssd1 vssd1 vccd1 vccd1 _0119_ sky130_fd_sc_hd__inv_2
XANTENNA__3362__B1 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2538_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0840_ _1235_ vssd1 vssd1
+ vccd1 vccd1 _0504_ sky130_fd_sc_hd__a21bo_1
X_4590__454 vssd1 vssd1 vccd1 vccd1 net454 _4590__454/LO sky130_fd_sc_hd__conb_1
X_4208_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[70\]
+ _0197_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[70\] sky130_fd_sc_hd__dfrtp_1
X_2469_ team_10_WB.instance_to_wrap.host_row1\[58\] net132 net128 team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\]
+ _1208_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__a221o_1
XANTENNA__4167__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4139_ clknet_leaf_9_wb_clk_i _0610_ _0138_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3353__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout181 _1709_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
Xfanout170 _1702_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_4
Xfanout192 _0994_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_4
XANTENNA__3997__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2459__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2919__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ net250 vssd1 vssd1 vccd1 vccd1 _0042_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4490_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[47\]
+ _0473_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_3441_ net181 _1802_ _1809_ net173 vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__a22o_1
XANTENNA__3344__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3372_ team_10_WB.instance_to_wrap.host_row2\[50\] net170 net179 team_10_WB.instance_to_wrap.host_row2\[66\]
+ _1749_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__a221o_1
X_2323_ _1097_ _1098_ _0868_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2254_ team_10_WB.instance_to_wrap.gamelogic.setWord\[35\] net215 vssd1 vssd1 vccd1
+ vccd1 _1036_ sky130_fd_sc_hd__nand2_1
XANTENNA__4002__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2185_ _0919_ _0972_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4152__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_62_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout232_A _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1969_ team_10_WB.instance_to_wrap.gamelogic.setWord\[18\] net147 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[26\]
+ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__o22a_1
XANTENNA__2386__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3708_ net235 vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_961 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4688_ net183 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout118_X net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3639_ net282 vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3102__A3 net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3326__B1 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4025__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 team_10_WB.instance_to_wrap.keypadFSMHost.strobe_edge vssd1 vssd1 vccd1 vccd1
+ net461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4175__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2301__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2266__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[27\]
+ _0058_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_2941_ net213 net154 net122 net661 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[46\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4611_ net386 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
X_2872_ net193 _1458_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[0\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__3097__B net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3014__C1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4270__Q team_10_WB.instance_to_wrap.gamelogic.letter\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4542_ net354 vssd1 vssd1 vccd1 vccd1 DAT_O[16] sky130_fd_sc_hd__buf_2
XFILLER_0_5_758 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4473_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[30\]
+ _0456_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3424_ team_10_WB.instance_to_wrap.host_row1\[77\] net302 _1708_ vssd1 vssd1 vccd1
+ vccd1 _1799_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3841__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3355_ team_10_WB.instance_to_wrap.dispFSM.guesses\[65\] _1719_ _1733_ net232 vssd1
+ vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__a211o_1
X_3286_ net295 _1670_ _1671_ vssd1 vssd1 vccd1 vccd1 _0567_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_55_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _0841_ _1073_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2237_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _0799_ _0805_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\]
+ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__a221o_1
XANTENNA__3052__S net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout182_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2168_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4672__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2099_ team_10_WB.instance_to_wrap.dispFSM.guesses\[21\] net143 net107 net562 vssd1
+ vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3020__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4048__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4198__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2047__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3140_ _0889_ _0894_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__or2_1
XANTENNA__2522__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3071_ team_10_WB.instance_to_wrap.gamelogic.setWord\[32\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2022_ _0892_ _0896_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_18_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3973_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[10\]
+ _0041_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_46_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2924_ net615 net156 net125 net625 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[29\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2855_ net708 _1447_ net176 vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4525_ net337 vssd1 vssd1 vccd1 vccd1 CYC_O sky130_fd_sc_hd__buf_2
XFILLER_0_53_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold201 team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] vssd1 vssd1 vccd1 vccd1
+ net658 sky130_fd_sc_hd__dlygate4sd3_1
X_2786_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\] vssd1 vssd1 vccd1 vccd1 _1396_
+ sky130_fd_sc_hd__or3_1
XANTENNA__2210__B1 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold223 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\] vssd1 vssd1 vccd1
+ vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold234 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\] vssd1 vssd1 vccd1
+ vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold212 team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] vssd1 vssd1 vccd1 vccd1
+ net669 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold245 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] vssd1 vssd1 vccd1 vccd1
+ net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] vssd1 vssd1 vccd1 vccd1
+ net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\] vssd1 vssd1 vccd1
+ vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ clknet_leaf_27_wb_clk_i net617 _0439_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold278 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\] vssd1 vssd1 vccd1
+ vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4340__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3407_ net67 net178 _1783_ net230 vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__o211a_1
X_4387_ clknet_leaf_6_wb_clk_i _0772_ _0370_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[24\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4667__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3338_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net211 _1707_ vssd1 vssd1
+ vccd1 vccd1 _1718_ sky130_fd_sc_hd__or3_2
XPHY_EDGE_ROW_37_Left_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4513__325 vssd1 vssd1 vccd1 vccd1 _4513__325/HI net325 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_5_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4490__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3269_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\]
+ _1657_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout185_X net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_764 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Left_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Left_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2268__B1 net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2825__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_wb_clk_i_X clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3420__S net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3480__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2440__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2991__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_2640_ _0926_ net189 vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__nand2_1
XANTENNA__4363__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2571_ team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] _0898_ vssd1 vssd1
+ vccd1 vccd1 _1256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4310_ clknet_leaf_17_wb_clk_i _0700_ _0299_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[33\]
+ sky130_fd_sc_hd__dfstp_1
X_4241_ clknet_leaf_30_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[5\]
+ _0230_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4172_ clknet_leaf_26_wb_clk_i _0641_ _0161_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3123_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] _1288_ _1553_ _0825_
+ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__o31a_1
X_3054_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] _1521_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[63\] sky130_fd_sc_hd__mux2_1
X_2005_ net221 net222 net223 vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__or3_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3471__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2454__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3956_ clknet_leaf_27_wb_clk_i _0007_ _0024_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_2907_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[20\] net153 net124 net691
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[12\]
+ sky130_fd_sc_hd__o22a_1
X_3887_ net277 vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__inv_2
XANTENNA__3566__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4658__427 vssd1 vssd1 vccd1 vccd1 _4658__427/HI net427 sky130_fd_sc_hd__conb_1
X_2838_ _1407_ _0515_ _1426_ _1409_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__o31a_1
X_2769_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[25\]
+ team_10_WB.instance_to_wrap.clock_div.count\[24\] _1380_ vssd1 vssd1 vccd1 vccd1
+ _1384_ sky130_fd_sc_hd__and4_1
X_4508_ net320 vssd1 vssd1 vccd1 vccd1 ADR_O[15] sky130_fd_sc_hd__buf_2
X_4439_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[36\]
+ _0422_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_38_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3462__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4386__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2489__B1 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3150__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3810_ net294 vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_29 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3741_ net285 vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_45_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2964__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3672_ net248 vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2623_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1074_ _1296_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0010_ sky130_fd_sc_hd__a22o_1
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[5] sky130_fd_sc_hd__buf_2
XFILLER_0_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4109__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2554_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] _1241_ vssd1 vssd1 vccd1
+ vccd1 _1246_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2485_ net540 net133 _1187_ _1215_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4224_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[86\]
+ _0213_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[86\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__4259__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4155_ clknet_leaf_28_wb_clk_i _0626_ _0145_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.strobe
+ sky130_fd_sc_hd__dfrtp_1
X_3106_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[11\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[12\]
+ _1546_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[13\] vssd1 vssd1 vccd1 vccd1
+ _1547_ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4086_ clknet_leaf_12_wb_clk_i _0557_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout262_A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3037_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__mux2_1
XANTENNA__3444__A2 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4680__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3939_ net237 vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4519__331 vssd1 vssd1 vccd1 vccd1 _4519__331/HI net331 sky130_fd_sc_hd__conb_1
XFILLER_0_30_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4363__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4606__381 vssd1 vssd1 vccd1 vccd1 _4606__381/HI net381 sky130_fd_sc_hd__conb_1
Xinput16 wbs_adr_i[17] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_1
Xinput27 wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_1
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3371__A1 team_10_WB.instance_to_wrap.host_row2\[82\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4401__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2270_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net213 vssd1 vssd1 vccd1
+ vccd1 _1052_ sky130_fd_sc_hd__or2_1
XANTENNA__2269__B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4583__451 vssd1 vssd1 vccd1 vccd1 net451 _4583__451/LO sky130_fd_sc_hd__conb_1
XANTENNA__1988__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4273__Q team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] net148 vssd1 vssd1 vccd1
+ vccd1 _0882_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2937__A1 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3724_ net244 vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3655_ net259 vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__inv_2
X_2606_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] _1287_ vssd1 vssd1
+ vccd1 vccd1 _1288_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3586_ net261 vssd1 vssd1 vccd1 vccd1 _0118_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3055__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2537_ _0871_ _1073_ _1088_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__nand3_1
X_2468_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] net197 vssd1 vssd1
+ vccd1 vccd1 _1208_ sky130_fd_sc_hd__and2_1
XANTENNA__3114__A1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4207_ clknet_leaf_25_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\]
+ _0196_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[69\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2399_ team_10_WB.instance_to_wrap.clock_div.count\[4\] team_10_WB.instance_to_wrap.clock_div.count\[6\]
+ team_10_WB.instance_to_wrap.clock_div.count\[5\] vssd1 vssd1 vccd1 vccd1 _1162_
+ sky130_fd_sc_hd__or3b_1
X_4138_ clknet_leaf_10_wb_clk_i _0609_ _0137_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3417__A2 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4069_ clknet_leaf_22_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[0\]
+ _0089_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__1979__A2 net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4424__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3754__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input38_A wbs_adr_i[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout171 _1702_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
Xfanout160 net164 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout193 _1222_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3408__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3041__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3440_ _1707_ _1804_ _1814_ _1717_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3371_ team_10_WB.instance_to_wrap.host_row2\[82\] net173 _1708_ team_10_WB.instance_to_wrap.host_row1\[74\]
+ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2322_ _0844_ _0851_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nand2_1
X_2253_ team_10_WB.instance_to_wrap.gamelogic.setWord\[36\] net214 vssd1 vssd1 vccd1
+ vccd1 _1035_ sky130_fd_sc_hd__xnor2_1
X_2184_ net134 _0972_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__and2_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4447__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1968_ team_10_WB.instance_to_wrap.gamelogic.setWord\[19\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[27\]
+ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4687_ net182 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_1
X_3707_ net235 vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1899_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\] vssd1 vssd1 vccd1 vccd1
+ _0823_ sky130_fd_sc_hd__inv_2
X_3638_ net280 vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3569_ net270 vssd1 vssd1 vccd1 vccd1 _0101_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3964__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] vssd1 vssd1 vccd1 vccd1 net462
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3659__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] net156 net125 net654 vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[45\] sky130_fd_sc_hd__a22o_1
XFILLER_0_29_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2871_ net1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[0\] _1457_ vssd1 vssd1 vccd1
+ vccd1 _1458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4610_ net385 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4541_ net353 vssd1 vssd1 vccd1 vccd1 DAT_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_29_Left_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_921 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4472_ clknet_leaf_27_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[29\]
+ _0455_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3423_ net68 net177 _1798_ net231 vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4619__391 vssd1 vssd1 vccd1 vccd1 _4619__391/HI net391 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_55_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] net173 _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3285_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[16\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\]
+ _1666_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2305_ _0841_ _0860_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nor2_1
X_2236_ _0796_ net212 net215 _0797_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__a22o_1
XANTENNA__3096__A3 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2167_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2098_ team_10_WB.instance_to_wrap.dispFSM.guesses\[14\] net112 net138 net579 vssd1
+ vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4626__395 vssd1 vssd1 vccd1 vccd1 _4626__395/HI net395 sky130_fd_sc_hd__conb_1
XFILLER_0_61_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout130_X net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_wb_clk_i_X clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3244__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_868 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4142__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3070_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _1529_ net202 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[71\] sky130_fd_sc_hd__mux2_1
X_2021_ _0892_ _0894_ net227 vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__or3b_1
XANTENNA__4292__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3972_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[9\]
+ _0040_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2923_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[36\] net152 net121 net681
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2854_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[5\]
+ _1444_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2785_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\]
+ _1394_ vssd1 vssd1 vccd1 vccd1 _1395_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4524_ net336 vssd1 vssd1 vccd1 vccd1 ADR_O[31] sky130_fd_sc_hd__buf_2
Xhold202 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[32\] vssd1 vssd1 vccd1
+ vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold213 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\] vssd1 vssd1 vccd1
+ vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold224 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\] vssd1 vssd1 vccd1
+ vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold235 team_10_WB.instance_to_wrap.dispFSM.guesses\[46\] vssd1 vssd1 vccd1 vccd1
+ net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4455_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[12\]
+ _0438_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\]
+ sky130_fd_sc_hd__dfstp_1
Xhold246 team_10_WB.instance_to_wrap.dispFSM.guesses\[68\] vssd1 vssd1 vccd1 vccd1
+ net703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\] vssd1 vssd1 vccd1 vccd1
+ net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] vssd1 vssd1 vccd1 vccd1
+ net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3406_ net232 _1774_ _1782_ _1767_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__a211o_1
X_4386_ clknet_leaf_1_wb_clk_i _0771_ _0369_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[23\]
+ sky130_fd_sc_hd__dfrtp_2
X_3337_ _1694_ _1714_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nor2_4
XFILLER_0_42_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2468__A team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4552__364 vssd1 vssd1 vccd1 vccd1 _4552__364/HI net364 sky130_fd_sc_hd__conb_1
XANTENNA__3063__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3268_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ net618 vssd1 vssd1
+ vccd1 vccd1 _1659_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2187__B net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout178_X net178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3199_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\] _1392_ vssd1 vssd1 vccd1
+ vccd1 _1617_ sky130_fd_sc_hd__xnor2_1
X_2219_ net28 net29 vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__nand2_1
XANTENNA__3474__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4015__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4165__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2201__A1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input20_A wbs_adr_i[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2268__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3937__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2955__A2_N _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_643 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4495__307 vssd1 vssd1 vccd1 vccd1 _4495__307/HI net307 sky130_fd_sc_hd__conb_1
XFILLER_0_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2570_ net223 net227 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[0\] vssd1
+ vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4536__348 vssd1 vssd1 vccd1 vccd1 _4536__348/HI net348 sky130_fd_sc_hd__conb_1
X_4240_ clknet_leaf_31_wb_clk_i team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[4\]
+ _0229_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.Rx_byte\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4171_ clknet_leaf_25_wb_clk_i _0640_ _0160_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\]
+ sky130_fd_sc_hd__dfstp_2
X_3122_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[1\] _1552_ _0824_ vssd1
+ vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_2_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4276__Q team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3456__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3053_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[23\]
+ net189 vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__mux2_1
X_2004_ net301 net3 vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__nand2_1
XANTENNA__4038__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3955_ clknet_leaf_27_wb_clk_i _0006_ _0023_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2906_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[19\] net153 net121 net724
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[11\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4188__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3886_ net263 vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2837_ _1407_ _1436_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2768_ team_10_WB.instance_to_wrap.clock_div.count\[24\] _1382_ net707 vssd1 vssd1
+ vccd1 vccd1 _1383_ sky130_fd_sc_hd__a21oi_1
X_4507_ net319 vssd1 vssd1 vccd1 vccd1 ADR_O[14] sky130_fd_sc_hd__buf_2
X_2699_ _0807_ team_10_WB.instance_to_wrap.message_reg.state\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ _1343_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _1344_ sky130_fd_sc_hd__o221a_1
X_4438_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[35\]
+ _0421_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4369_ clknet_leaf_26_wb_clk_i _0754_ _0352_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\]
+ sky130_fd_sc_hd__dfstp_2
XPHY_EDGE_ROW_16_Left_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3447__B1 net168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2645__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4641__410 vssd1 vssd1 vccd1 vccd1 _4641__410/HI net410 sky130_fd_sc_hd__conb_1
XFILLER_0_64_576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2489__B2 team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4330__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_19 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3740_ net286 vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3671_ net258 vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4480__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2622_ _1116_ _1235_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nor2_1
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[6] sky130_fd_sc_hd__buf_2
XFILLER_0_2_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2553_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2484_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\] _0991_ vssd1 vssd1 vccd1
+ vccd1 _1215_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4223_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\]
+ _0212_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[85\] sky130_fd_sc_hd__dfrtp_1
X_4154_ clknet_leaf_11_wb_clk_i _0625_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfxtp_1
X_4085_ clknet_leaf_12_wb_clk_i _0556_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3105_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1396_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[10\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\]
+ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__o2111a_1
X_3036_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] _1512_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[54\] sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2465__B net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3938_ net242 vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3869_ net261 vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4558__370 vssd1 vssd1 vccd1 vccd1 _4558__370/HI net370 sky130_fd_sc_hd__conb_1
XANTENNA__4203__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__2891__A1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Left_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3487__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 wbs_adr_i[28] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_1
Xinput17 wbs_adr_i[18] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput39 wbs_adr_i[9] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_793 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_16 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3426__S net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3371__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3014__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1984_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] net149 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\]
+ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__o22a_1
X_3723_ net244 vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3654_ net256 vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__inv_2
XANTENNA__4226__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2605_ _0888_ _1279_ _0900_ _0899_ _0895_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_11_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3585_ net280 vssd1 vssd1 vccd1 vccd1 _0117_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3362__A2 net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2536_ net479 team_10_WB.instance_to_wrap.buffer.temp_guess\[0\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0505_ sky130_fd_sc_hd__mux2_1
X_2467_ net555 net129 _1207_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__o21a_1
X_4206_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[68\]
+ _0195_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[68\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__4376__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2398_ team_10_WB.instance_to_wrap.clock_div.count\[8\] team_10_WB.instance_to_wrap.clock_div.count\[13\]
+ team_10_WB.instance_to_wrap.clock_div.count\[12\] vssd1 vssd1 vccd1 vccd1 _1161_
+ sky130_fd_sc_hd__or3_1
X_4137_ clknet_leaf_7_wb_clk_i _0608_ _0136_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4068_ clknet_leaf_31_wb_clk_i _0550_ _0088_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3019_ team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] net190 vssd1 vssd1 vccd1
+ vccd1 _1504_ sky130_fd_sc_hd__or2_1
XANTENNA__4691__A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4226__439 vssd1 vssd1 vccd1 vccd1 net439 _4226__439/LO sky130_fd_sc_hd__conb_1
XFILLER_0_61_343 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3353__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2561__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 _1612_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
Xfanout161 net163 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout183 net184 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout150 _0862_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout194 _0991_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__buf_4
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3344__A2 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ team_10_WB.instance_to_wrap.host_row1\[42\] _1693_ net174 team_10_WB.instance_to_wrap.host_row2\[42\]
+ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2321_ _0819_ _0849_ _0851_ _0867_ vssd1 vssd1 vccd1 vccd1 _1097_ sky130_fd_sc_hd__or4_1
X_2252_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] _1033_ _1025_ _1027_
+ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2183_ _0923_ _0947_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1967_ team_10_WB.instance_to_wrap.gamelogic.setWord\[20\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[28\]
+ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout120_A net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ net239 vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__inv_2
X_4686_ net183 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_1
X_1898_ net219 vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3637_ net256 vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__inv_2
XANTENNA__3066__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3568_ net270 vssd1 vssd1 vccd1 vccd1 _0100_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4686__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2519_ net543 _1231_ _1232_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] vssd1 vssd1
+ vccd1 vccd1 _0526_ sky130_fd_sc_hd__a22o_1
X_3499_ net251 vssd1 vssd1 vccd1 vccd1 _0031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_30_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3326__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4369__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold6 _0511_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4071__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2870_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ net224 vssd1 vssd1 vccd1 vccd1 _1457_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540_ net352 vssd1 vssd1 vccd1 vccd1 DAT_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_40_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4471_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[28\]
+ _0454_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3422_ net232 _1788_ _1794_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3353_ team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] net180 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[9\]
+ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3284_ net702 _1668_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _0868_ _1080_ _1081_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2235_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _0800_ _0803_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1017_ sky130_fd_sc_hd__a22o_1
X_2166_ _0936_ _0939_ _0954_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__a21o_1
XANTENNA__4414__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2097_ team_10_WB.instance_to_wrap.dispFSM.guesses\[23\] net145 net108 net577 vssd1
+ vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2461__C1 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2999_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\] net165 _1497_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[32\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3005__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4669_ net432 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_4_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4189__Q team_10_WB.instance_to_wrap.host_row2\[51\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4094__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_wb_clk_i_X clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_30_Left_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3434__S net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4437__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2020_ _0899_ _0902_ _0901_ _0896_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__and4bb_4
XTAP_TAPCELL_ROW_50_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3971_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[8\]
+ _0039_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_2922_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\] net151 net120 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[27\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2853_ _1447_ net176 _1446_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[4\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2784_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ vssd1 vssd1 vccd1 vccd1 _1394_ sky130_fd_sc_hd__or4_1
X_4523_ net335 vssd1 vssd1 vccd1 vccd1 ADR_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold225 team_10_WB.instance_to_wrap.dispFSM.guesses\[20\] vssd1 vssd1 vccd1 vccd1
+ net682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold203 team_10_WB.instance_to_wrap.dispFSM.guesses\[9\] vssd1 vssd1 vccd1 vccd1
+ net660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 team_10_WB.instance_to_wrap.dispFSM.guesses\[14\] vssd1 vssd1 vccd1 vccd1
+ net671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold269 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[9\] vssd1 vssd1 vccd1 vccd1
+ net726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 team_10_WB.instance_to_wrap.dispFSM.guesses\[8\] vssd1 vssd1 vccd1 vccd1
+ net704 sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[11\]
+ _0437_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[11\]
+ sky130_fd_sc_hd__dfstp_1
Xhold258 team_10_WB.instance_to_wrap.dispFSM.guesses\[49\] vssd1 vssd1 vccd1 vccd1
+ net715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] vssd1 vssd1 vccd1
+ vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
X_4385_ clknet_leaf_7_wb_clk_i _0770_ _0368_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\]
+ sky130_fd_sc_hd__dfstp_2
X_3405_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\] _1690_ net175 _1775_
+ _1781_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkload22_A clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3336_ team_10_WB.instance_to_wrap.dispFSM.guesses\[48\] net167 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[72\]
+ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a22o_1
XANTENNA__2468__B net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3267_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ _1658_ vssd1 vssd1
+ vccd1 vccd1 _0561_ sky130_fd_sc_hd__o21a_1
X_3198_ _1393_ _1611_ _1616_ vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__and3_1
X_2218_ net25 net24 net27 net26 vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2149_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] _0943_ vssd1 vssd1 vccd1
+ vccd1 _0944_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3954__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1960__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1960__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2268__A2 _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3465__A1 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input13_A wbs_adr_i[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4170_ clknet_leaf_25_wb_clk_i _0639_ _0159_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_TAPCELL_ROW_52_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3121_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\] _1860_ vssd1 vssd1
+ vccd1 vccd1 _1552_ sky130_fd_sc_hd__and2b_1
XANTENNA__2900__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3052_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] _1520_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[62\] sky130_fd_sc_hd__mux2_1
XANTENNA__3977__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1920__B net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2003_ team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_26_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3954_ clknet_leaf_25_wb_clk_i _0005_ _0022_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.state\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_2905_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[18\] net153 net121 net697
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[10\]
+ sky130_fd_sc_hd__o22a_1
X_3885_ net269 vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__inv_2
X_2836_ _1436_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2767_ net603 _1382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[24\]
+ sky130_fd_sc_hd__xor2_1
X_4506_ net318 vssd1 vssd1 vccd1 vccd1 ADR_O[13] sky130_fd_sc_hd__buf_2
XANTENNA__3392__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout200_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2698_ team_10_WB.instance_to_wrap.message_reg.msg\[0\] team_10_WB.instance_to_wrap.message_reg.msg\[1\]
+ team_10_WB.instance_to_wrap.message_reg.msg\[2\] team_10_WB.instance_to_wrap.message_reg.msg\[3\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__mux4_1
X_4437_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[34\]
+ _0420_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input5_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4368_ clknet_leaf_26_wb_clk_i _0753_ _0351_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_3319_ _1688_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout190_X net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4299_ clknet_leaf_20_wb_clk_i _0689_ _0288_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2645__C team_10_WB.instance_to_wrap.host_message_reg.Cstate vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4132__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4282__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1050 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2587__A1_N net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4377__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2489__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3438__A1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input16_X net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3438__B2 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2949__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4503__315 vssd1 vssd1 vccd1 vccd1 _4503__315/HI net315 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_45_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3670_ net241 vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3683__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2621_ _0006_ _0009_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMHost.next_state\[2\]
+ sky130_fd_sc_hd__or2_1
XFILLER_0_24_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_3_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2552_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\] _1243_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__a21o_1
X_4222_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[84\]
+ _0211_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[84\] sky130_fd_sc_hd__dfrtp_1
X_2483_ net535 net130 _1185_ _1214_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__a22o_1
X_4153_ clknet_leaf_11_wb_clk_i _0624_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ clknet_leaf_14_wb_clk_i _0555_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_3104_ team_10_WB.EN_VAL_REG net182 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__or2_1
XANTENNA__3429__A1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3035_ team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4155__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3937_ net241 vssd1 vssd1 vccd1 vccd1 _0469_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout248_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3069__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3868_ net275 vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2819_ _1421_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3799_ net281 vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__inv_2
XANTENNA__4689__A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input8_X net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 wbs_adr_i[19] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4028__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4178__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4648__417 vssd1 vssd1 vccd1 vccd1 _4648__417/HI net417 sky130_fd_sc_hd__conb_1
XFILLER_0_59_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1983_ team_10_WB.instance_to_wrap.gamelogic.setWord\[15\] _0874_ _0881_ net159 vssd1
+ vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__o211a_1
X_3722_ net244 vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3653_ net256 vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2604_ _1268_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[0\] _1265_ vssd1
+ vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_11_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3584_ net262 vssd1 vssd1 vccd1 vccd1 _0116_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2535_ net476 team_10_WB.instance_to_wrap.buffer.temp_guess\[1\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0506_ sky130_fd_sc_hd__mux2_1
X_2466_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] net197 _1187_
+ _1206_ net132 vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4205_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[67\]
+ _0194_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[67\] sky130_fd_sc_hd__dfrtp_1
X_4136_ clknet_leaf_2_wb_clk_i _0607_ _0135_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_2397_ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[2\]
+ team_10_WB.instance_to_wrap.clock_div.count\[9\] team_10_WB.instance_to_wrap.clock_div.count\[10\]
+ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__or4bb_1
XANTENNA__2476__B net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4067_ clknet_leaf_31_wb_clk_i _0549_ _0087_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_3018_ net197 _1503_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[45\]
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout153_X net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout173 _1701_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_4
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
Xfanout151 net153 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
Xfanout184 net101 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__clkbuf_8
Xfanout195 _0885_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_2
XFILLER_0_9_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3498__A net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4006__RESET_B net274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2001__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2320_ _1094_ _1095_ _0869_ _1092_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__o2bb2a_1
X_2251_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] _0798_ _0800_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\]
+ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2182_ team_10_WB.instance_to_wrap.gamelogic.state\[0\] net218 team_10_WB.instance_to_wrap.gamelogic.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4509__321 vssd1 vssd1 vccd1 vccd1 _4509__321/HI net321 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_62_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1966_ team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] _0874_ _0878_ net157 vssd1
+ vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3705_ net239 vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4685_ net437 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_0_43_355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1897_ net300 vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__inv_2
X_3636_ net277 vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3567_ net290 vssd1 vssd1 vccd1 vccd1 _0099_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2518_ _0807_ _0808_ net145 vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__and3_2
X_3498_ net290 vssd1 vssd1 vccd1 vccd1 _0030_ sky130_fd_sc_hd__inv_2
X_2449_ net572 net132 _1191_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ _1190_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__a221o_1
XANTENNA__3082__S net202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4119_ clknet_leaf_8_wb_clk_i _0590_ _0118_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3008__C1 net206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A wbs_we_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4385__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 team_10_WB.instance_to_wrap.clock_div.count\[29\] vssd1 vssd1 vccd1 vccd1 net464
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4216__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4366__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3014__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4470_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[27\]
+ _0453_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3421_ net179 _1795_ _1796_ net175 _1781_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3352_ team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] net174 _1715_ team_10_WB.instance_to_wrap.dispFSM.guesses\[73\]
+ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2525__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[1\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2303_ net225 net226 _0869_ vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__or3_1
X_3283_ net517 _1666_ _1669_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_55_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] _0805_ vssd1 vssd1 vccd1
+ vccd1 _1016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2165_ _0942_ _0955_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 _0656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2096_ team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] net114 net141 net727 vssd1
+ vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout230_A _0018_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3866__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2998_ net126 _1496_ vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__nand2_2
XANTENNA__3077__S net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1949_ _0841_ _0871_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__nor2_1
X_4668_ net184 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3619_ net269 vssd1 vssd1 vccd1 vccd1 _0151_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4599_ net199 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_1
XANTENNA__3477__C1 net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2945__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4389__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_336 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1963__C1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3483__A2 _1853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3970_ clknet_leaf_28_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[7\]
+ _0038_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2921_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\] net151 net120 net709
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[26\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_31 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2852_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[3\]
+ _1442_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__and3_1
X_2783_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4522_ net334 vssd1 vssd1 vccd1 vccd1 ADR_O[29] sky130_fd_sc_hd__buf_2
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold204 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] vssd1 vssd1 vccd1
+ vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold226 team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] vssd1 vssd1 vccd1 vccd1
+ net683 sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[10\]
+ _0436_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[10\]
+ sky130_fd_sc_hd__dfstp_1
Xhold215 team_10_WB.instance_to_wrap.dispFSM.guesses\[78\] vssd1 vssd1 vccd1 vccd1
+ net672 sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _1777_ _1780_ net177 vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__o21ai_2
Xhold237 team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] vssd1 vssd1 vccd1 vccd1
+ net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] vssd1 vssd1 vccd1 vccd1
+ net705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold259 team_10_WB.instance_to_wrap.clock_div.count\[14\] vssd1 vssd1 vccd1 vccd1
+ net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4384_ clknet_leaf_27_wb_clk_i _0769_ _0367_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_892 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload15_A clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3335_ _1687_ _1714_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__nor2_4
X_3266_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[10\] _1657_ net296 vssd1 vssd1
+ vccd1 vccd1 _1658_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2217_ net15 net17 net18 net16 vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__or4bb_1
X_3197_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1616_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3474__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2484__B _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2148_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__nand2_1
X_2079_ team_10_WB.instance_to_wrap.dispFSM.guesses\[33\] net109 net135 team_10_WB.instance_to_wrap.dispFSM.guesses\[41\]
+ vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_984 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4061__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2976__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_951 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4404__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3120_ net195 _1550_ _1290_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__o21ba_1
X_3051_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[22\]
+ net190 vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__mux2_1
XANTENNA__3456__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2002_ team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge1 team_10_WB.instance_to_wrap.keypadFSMPlayer.strobe_edge
+ vssd1 vssd1 vccd1 vccd1 _0885_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3953_ clknet_leaf_23_wb_clk_i _0016_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2904_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\] net154 net122 net670
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[9\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3884_ net275 vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__inv_2
X_2835_ _1415_ _1426_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4084__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2766_ _1381_ _1382_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[23\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4505_ net317 vssd1 vssd1 vccd1 vccd1 ADR_O[12] sky130_fd_sc_hd__buf_2
XFILLER_0_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2697_ _1341_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[2\] vssd1 vssd1
+ vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2b_1
X_4436_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[33\]
+ _0419_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4367_ clknet_leaf_2_wb_clk_i _0752_ _0350_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[4\]
+ sky130_fd_sc_hd__dfstp_1
X_3318_ _1697_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4298_ clknet_leaf_19_wb_clk_i net598 _0287_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3249_ _1610_ _1647_ net298 vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2495__A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3447__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4427__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3383__A1 net303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3383__B2 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4393__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3013__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2949__B2 net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4542__354 vssd1 vssd1 vccd1 vccd1 _4542__354/HI net354 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_45_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2620_ _0840_ _0860_ _1295_ _1085_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[4\]
+ vssd1 vssd1 vccd1 vccd1 _0009_ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2551_ _1239_ _1242_ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_50_294 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2482_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] net186 vssd1 vssd1 vccd1
+ vccd1 _1214_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4221_ clknet_leaf_5_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[83\]
+ _0210_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[83\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3944__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ clknet_leaf_11_wb_clk_i _0623_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__dfxtp_1
X_4083_ clknet_leaf_13_wb_clk_i _0554_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__3429__A2 team_10_WB.instance_to_wrap.host_row2\[101\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_3103_ net157 _1302_ net198 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_state
+ sky130_fd_sc_hd__mux2_1
X_3034_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] _1511_ net208 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[53\] sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2101__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3936_ net240 vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout143_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3867_ net261 vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3874__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2818_ _1410_ _1422_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__nand2_1
X_3798_ net294 vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2749_ team_10_WB.instance_to_wrap.clock_div.count\[18\] _1370_ vssd1 vssd1 vccd1
+ vccd1 _1371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_X clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3085__S net189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3117__A1 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4419_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[16\]
+ _0402_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4526__338 vssd1 vssd1 vccd1 vccd1 _4526__338/HI net338 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_24_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_25_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput19 wbs_adr_i[1] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3967__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4388__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1982_ team_10_WB.instance_to_wrap.gamelogic.setWord\[7\] net148 vssd1 vssd1 vccd1
+ vccd1 _0881_ sky130_fd_sc_hd__or2_1
X_3721_ net244 vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__inv_2
XANTENNA__3694__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3652_ net277 vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3583_ net276 vssd1 vssd1 vccd1 vccd1 _0115_ sky130_fd_sc_hd__inv_2
X_2603_ _0016_ _0013_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.next_state\[1\]
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2534_ net481 team_10_WB.instance_to_wrap.buffer.temp_guess\[2\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2465_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] net194 vssd1 vssd1 vccd1
+ vccd1 _1206_ sky130_fd_sc_hd__or2_1
XANTENNA__4122__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4631__400 vssd1 vssd1 vccd1 vccd1 _4631__400/HI net400 sky130_fd_sc_hd__conb_1
X_4204_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[66\]
+ _0193_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[66\] sky130_fd_sc_hd__dfrtp_1
X_2396_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _0854_ _1158_ net567 vssd1
+ vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__a22o_1
X_4135_ clknet_leaf_10_wb_clk_i _0606_ _0134_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ clknet_leaf_30_wb_clk_i _0548_ _0086_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout260_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3017_ team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[5\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3035__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3919_ net278 vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2013__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout152 net153 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout174 _1696_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_4
Xfanout141 net142 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout163 net164 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout185 _0995_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
Xfanout196 _0855_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3026__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3019__A team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4145__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2001__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2001__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2250_ team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] _0804_ _1029_ _1031_ vssd1
+ vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__a211o_1
XANTENNA__4295__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2181_ _0970_ team_10_WB.instance_to_wrap.correct\[0\] _0958_ vssd1 vssd1 vccd1 vccd1
+ _0653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4548__360 vssd1 vssd1 vccd1 vccd1 _4548__360/HI net360 sky130_fd_sc_hd__conb_1
XANTENNA__3017__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1965_ team_10_WB.instance_to_wrap.gamelogic.setWord\[21\] net147 vssd1 vssd1 vccd1
+ vccd1 _0878_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3704_ net235 vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__inv_2
XANTENNA__2532__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4684_ net182 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1896_ team_10_WB.instance_to_wrap.host_col\[0\] vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__inv_2
X_3635_ net264 vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3566_ net290 vssd1 vssd1 vccd1 vccd1 _0098_ sky130_fd_sc_hd__inv_2
X_2517_ team_10_WB.instance_to_wrap.message_reg.state\[1\] net145 _0808_ vssd1 vssd1
+ vccd1 vccd1 _1231_ sky130_fd_sc_hd__o21ai_4
X_3497_ net290 vssd1 vssd1 vccd1 vccd1 _0029_ sky130_fd_sc_hd__inv_2
X_2448_ net564 net130 _1187_ _1197_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__a22o_1
X_2379_ _1099_ _1151_ _1135_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__mux2_1
X_4118_ clknet_leaf_17_wb_clk_i _0589_ _0117_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[53\]
+ sky130_fd_sc_hd__dfrtp_1
X_4049_ clknet_leaf_14_wb_clk_i _0534_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4168__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1990__B1 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input36_A wbs_adr_i[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 team_10_WB.instance_to_wrap.buffer.Rx_byte\[7\] vssd1 vssd1 vccd1 vccd1 net465
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3247__B1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3021__B net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2470__B2 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2470__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2205__X _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1981__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3420_ team_10_WB.instance_to_wrap.host_row2\[44\] team_10_WB.instance_to_wrap.dispFSM.guesses\[20\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__mux2_1
X_3351_ net717 net178 _1730_ net231 vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_59_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2302_ _0844_ _0847_ _0853_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__o21a_1
X_3282_ net295 _1668_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_55_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _0797_ net215 _0804_ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] _1014_
+ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2164_ _0942_ _0943_ _0957_ _0955_ net675 vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__a32o_1
XFILLER_0_49_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2095_ team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] net110 net135 net700 vssd1
+ vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4310__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2461__B2 _1189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2997_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] _1494_ _1495_ vssd1
+ vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3410__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1948_ _0865_ _0870_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_17_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4460__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4667_ net184 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_1
X_1879_ net217 vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3618_ net251 vssd1 vssd1 vccd1 vccd1 _0150_ sky130_fd_sc_hd__inv_2
X_4598_ net199 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_1
X_3549_ net286 vssd1 vssd1 vccd1 vccd1 _0081_ sky130_fd_sc_hd__inv_2
XANTENNA__3477__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2945__B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4396__Q team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4333__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2920_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[33\] net154 net123 net665
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[25\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4483__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_43 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2851_ team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[4\] _1444_ vssd1 vssd1
+ vccd1 vccd1 _1446_ sky130_fd_sc_hd__or2_1
X_2782_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\] _1391_ vssd1 vssd1 vccd1
+ vccd1 _1392_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ net333 vssd1 vssd1 vccd1 vccd1 ADR_O[28] sky130_fd_sc_hd__buf_2
X_4452_ clknet_leaf_11_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[9\]
+ _0435_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[9\]
+ sky130_fd_sc_hd__dfstp_1
Xhold216 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[35\] vssd1 vssd1 vccd1
+ vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 team_10_WB.instance_to_wrap.dispFSM.guesses\[17\] vssd1 vssd1 vccd1 vccd1
+ net662 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold249 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ net706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 team_10_WB.instance_to_wrap.dispFSM.guesses\[16\] vssd1 vssd1 vccd1 vccd1
+ net695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 team_10_WB.instance_to_wrap.dispFSM.guesses\[72\] vssd1 vssd1 vccd1 vccd1
+ net684 sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _1685_ _1720_ _1778_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__or4_1
X_4383_ clknet_leaf_6_wb_clk_i _0768_ _0366_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[20\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3334_ _1707_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] net210 vssd1 vssd1
+ vccd1 vccd1 _1714_ sky130_fd_sc_hd__or3b_2
XFILLER_0_42_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3265_ net296 _1656_ _1657_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nor3_1
XANTENNA__3459__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2216_ net21 net20 net23 net22 vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__or4_1
X_3196_ _1391_ _1611_ _1615_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__and3b_1
XANTENNA_fanout173_A _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2147_ _0937_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__nor2_4
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2078_ team_10_WB.instance_to_wrap.dispFSM.guesses\[34\] net114 net141 net636 vssd1
+ vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4206__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4356__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_749 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output67_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2900__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3050_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] _1519_ net208 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[61\] sky130_fd_sc_hd__mux2_1
X_2001_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] net148 net118
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1 vccd1 _0748_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2805__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3952_ clknet_leaf_21_wb_clk_i _0015_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_2903_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[16\] net153 net124 net734
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[8\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3883_ net267 vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__inv_2
X_2834_ _0515_ _1428_ _1435_ _1411_ vssd1 vssd1 vccd1 vccd1 _0002_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_835 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_771 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4504_ net316 vssd1 vssd1 vccd1 vccd1 ADR_O[11] sky130_fd_sc_hd__buf_2
XFILLER_0_53_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_wb_clk_i_X clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2765_ team_10_WB.instance_to_wrap.clock_div.count\[23\] team_10_WB.instance_to_wrap.clock_div.count\[22\]
+ _1378_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__and3_1
XANTENNA__3392__A2 _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2696_ team_10_WB.instance_to_wrap.message_reg.msg\[4\] team_10_WB.instance_to_wrap.message_reg.msg\[5\]
+ team_10_WB.instance_to_wrap.message_reg.msg\[6\] team_10_WB.instance_to_wrap.message_reg.msg\[7\]
+ team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[0\] team_10_WB.instance_to_wrap.uart_transmitter.bit_index\[1\]
+ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__mux4_1
X_4435_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[32\]
+ _0418_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4379__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4366_ clknet_leaf_2_wb_clk_i _0751_ _0349_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3317_ _0815_ net211 _1680_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__or3_2
XFILLER_0_6_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1951__Y _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4297_ clknet_leaf_12_wb_clk_i _0687_ _0286_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[20\]
+ sky130_fd_sc_hd__dfstp_1
X_3248_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[3\] _1608_ vssd1 vssd1 vccd1
+ vccd1 _1647_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2495__B _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3179_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] _1602_ vssd1 vssd1 vccd1 vccd1
+ _0503_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2016__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3368__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2550_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2481_ net551 net133 _1187_ _1213_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__a22o_1
X_4220_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[82\]
+ _0209_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[82\] sky130_fd_sc_hd__dfrtp_1
X_4151_ clknet_leaf_11_wb_clk_i _0622_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__dfxtp_1
X_4082_ clknet_leaf_13_wb_clk_i _0553_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3102_ net202 net602 net189 _1545_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[87\]
+ sky130_fd_sc_hd__a31o_1
X_3033_ team_10_WB.instance_to_wrap.gamelogic.setWord\[13\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\]
+ net192 vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Left_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2535__S _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3935_ net277 vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__inv_2
XANTENNA__4051__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3866_ net265 vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout136_A net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2817_ _0516_ _1409_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3797_ net285 vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_52_Left_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2748_ _1369_ _1370_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[17\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4418_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[15\]
+ _0401_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_2679_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] _1327_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a21o_1
Xfanout301 net304 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_4
X_4349_ clknet_leaf_16_wb_clk_i _0739_ _0338_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[72\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2793__X _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__A2 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2564__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[3\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4074__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1981_ team_10_WB.instance_to_wrap.gamelogic.setWord\[8\] net150 net117 team_10_WB.instance_to_wrap.gamelogic.setWord\[16\]
+ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3720_ net244 vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3651_ net258 vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
X_3582_ net262 vssd1 vssd1 vccd1 vccd1 _0114_ sky130_fd_sc_hd__inv_2
X_2602_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\] _1275_ _1285_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ vssd1 vssd1 vccd1 vccd1 _0013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2533_ net470 team_10_WB.instance_to_wrap.buffer.temp_guess\[3\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2464_ net614 net129 _1194_ _1205_ vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__o22a_1
X_4203_ clknet_leaf_10_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[65\]
+ _0192_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[65\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2395_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked net226 _0850_ _1158_ net588
+ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__a32o_1
X_4134_ clknet_leaf_17_wb_clk_i _0605_ _0133_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4417__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ clknet_leaf_21_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[2\]
+ _0085_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3016_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[4\] net185 _1502_ net206
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\] sky130_fd_sc_hd__o211a_1
XANTENNA_fanout253_A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3885__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3918_ net243 vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3849_ net241 vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2013__B net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout131 _1183_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_4
Xfanout120 net121 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4097__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout153 _1182_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_4
Xfanout164 net166 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_2
Xfanout142 _0914_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
Xfanout175 _1696_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__buf_2
Xfanout186 _0995_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_2
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3019__B net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4654__423 vssd1 vssd1 vccd1 vccd1 _4654__423/HI net423 sky130_fd_sc_hd__conb_1
X_2180_ _0936_ _0961_ _0969_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2473__C1 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1964_ team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] net149 net118 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\]
+ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4683_ net436 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_50_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3703_ net235 vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1895_ team_10_WB.instance_to_wrap.host_col\[1\] vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3634_ net253 vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3565_ net290 vssd1 vssd1 vccd1 vccd1 _0097_ sky130_fd_sc_hd__inv_2
XANTENNA__1953__A net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2516_ net224 _1225_ _1230_ vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__a21oi_1
X_3496_ net290 vssd1 vssd1 vccd1 vccd1 _0028_ sky130_fd_sc_hd__inv_2
X_2447_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] net194 vssd1 vssd1 vccd1
+ vccd1 _1197_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2378_ _1130_ _1150_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__nor2_1
X_4117_ clknet_leaf_8_wb_clk_i _0588_ _0116_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_4048_ clknet_leaf_14_wb_clk_i _0533_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3957__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4638__407 vssd1 vssd1 vccd1 vccd1 _4638__407/HI net407 sky130_fd_sc_hd__conb_1
XFILLER_0_62_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1990__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1990__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2959__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4012__Q team_10_WB.instance_to_wrap.dispFSM.msg\[4\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold9 _0512_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input29_A wbs_adr_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2470__A2 net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4112__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4262__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3350_ _1726_ _1729_ net178 vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__or3b_1
XANTENNA__2930__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2301_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[6\] _1078_ _1076_
+ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__o21a_1
X_3281_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[14\]
+ _1664_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_55_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net214 vssd1 vssd1 vccd1
+ vccd1 _1014_ sky130_fd_sc_hd__xnor2_1
XANTENNA__2808__S _1403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2163_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__or2_1
X_2094_ team_10_WB.instance_to_wrap.dispFSM.guesses\[18\] net114 net142 net699 vssd1
+ vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_30 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2461__A2 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2996_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\] _0838_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[38\]
+ _0839_ net165 vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__a41o_1
XFILLER_0_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1947_ net2 net229 _0858_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__nor3_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4666_ net184 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_1
X_1878_ net216 vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout216_A team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4597_ net200 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_1
X_3617_ net269 vssd1 vssd1 vccd1 vccd1 _0149_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3548_ net286 vssd1 vssd1 vccd1 vccd1 _0080_ sky130_fd_sc_hd__inv_2
XANTENNA__2921__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3479_ team_10_WB.instance_to_wrap.host_row2\[79\] net167 _1849_ _1851_ vssd1 vssd1
+ vccd1 vccd1 _1852_ sky130_fd_sc_hd__a211o_1
XANTENNA__4135__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4285__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2204__A2 net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2850_ _1444_ _1445_ net176 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_clk_count\[3\]
+ sky130_fd_sc_hd__and3b_1
X_2781_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1391_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4520_ net332 vssd1 vssd1 vccd1 vccd1 ADR_O[27] sky130_fd_sc_hd__buf_2
XFILLER_0_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4451_ clknet_leaf_6_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[8\]
+ _0434_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[8\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__1954__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1954__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold217 team_10_WB.instance_to_wrap.dispFSM.guesses\[76\] vssd1 vssd1 vccd1 vccd1
+ net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] vssd1 vssd1 vccd1 vccd1
+ net663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] vssd1 vssd1 vccd1
+ vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\] _0815_ net211 _1690_
+ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__a31o_1
Xhold228 team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] vssd1 vssd1 vccd1 vccd1
+ net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2903__B1 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4382_ clknet_leaf_8_wb_clk_i _0767_ _0365_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[19\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4008__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3333_ team_10_WB.instance_to_wrap.host_row1\[40\] _1693_ _1700_ _1712_ vssd1 vssd1
+ vccd1 vccd1 _1713_ sky130_fd_sc_hd__a211o_2
XFILLER_0_0_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3264_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[9\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\]
+ _1653_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2215_ _0997_ _0998_ _0999_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__or4_2
XANTENNA__4158__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3195_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\] _1390_ vssd1 vssd1 vccd1
+ vccd1 _1615_ sky130_fd_sc_hd__or2_1
X_2146_ team_10_WB.instance_to_wrap.gamelogic.rights\[2\] _0939_ _0940_ vssd1 vssd1
+ vccd1 vccd1 _0941_ sky130_fd_sc_hd__or3_2
X_2077_ team_10_WB.instance_to_wrap.dispFSM.guesses\[35\] net112 net140 net646 vssd1
+ vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2979_ _0800_ _1488_ net158 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[21\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3395__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout121_X net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4649_ net418 vssd1 vssd1 vccd1 vccd1 la_data_out[19] sky130_fd_sc_hd__buf_2
XFILLER_0_13_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4570__446 vssd1 vssd1 vccd1 vccd1 net446 _4570__446/LO sky130_fd_sc_hd__conb_1
XANTENNA__2370__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_34_Left_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3386__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_463 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4300__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2000_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[1\] net148 net118
+ team_10_WB.instance_to_wrap.gamelogic.setWord\[1\] vssd1 vssd1 vccd1 vccd1 _0749_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__4450__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3951_ clknet_leaf_23_wb_clk_i _0014_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2902_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[15\] _1181_ net125 net501
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3882_ net275 vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2833_ _1423_ _1428_ _0518_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3377__B1 net179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2764_ team_10_WB.instance_to_wrap.clock_div.count\[23\] _1380_ vssd1 vssd1 vccd1
+ vccd1 _1381_ sky130_fd_sc_hd__nor2_1
X_4503_ net315 vssd1 vssd1 vccd1 vccd1 ADR_O[10] sky130_fd_sc_hd__buf_2
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2695_ _1239_ _1246_ _1010_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[2\]
+ sky130_fd_sc_hd__a21bo_1
X_4434_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[31\]
+ _0417_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4365_ clknet_leaf_1_wb_clk_i _0750_ _0348_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_3316_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4296_ clknet_leaf_16_wb_clk_i _0686_ _0285_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_3247_ _1610_ _1646_ net298 vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout283_A net299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_X clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3178_ _1277_ _1550_ _1551_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__o21ai_1
X_2129_ _0919_ _0929_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout169_X net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4473__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input11_A wbs_adr_i[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2207__A net194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3359__B1 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2480_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] net194 vssd1 vssd1 vccd1
+ vccd1 _1213_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4150_ clknet_leaf_11_wb_clk_i _0621_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__dfxtp_1
XANTENNA__3325__X _1705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[18] sky130_fd_sc_hd__clkbuf_4
X_3101_ _0788_ net202 vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__nor2_1
X_4081_ clknet_leaf_13_wb_clk_i _0552_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3032_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] _1510_ net205 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[52\] sky130_fd_sc_hd__mux2_1
XFILLER_0_53_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ net243 vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3865_ net275 vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2816_ _1416_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4346__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3796_ net286 vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout129_A _1184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3944__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ team_10_WB.instance_to_wrap.clock_div.count\[17\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ _1365_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2678_ net519 _1327_ _1330_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[6\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[14\]
+ _0400_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout302 net304 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input3_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4348_ clknet_leaf_19_wb_clk_i _0738_ _0337_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_4279_ clknet_leaf_15_wb_clk_i _0669_ _0268_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2645__A_N net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4219__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1980_ team_10_WB.instance_to_wrap.gamelogic.setWord\[9\] net149 net119 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\]
+ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__o22a_1
XANTENNA__4369__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2246__A1_N team_10_WB.instance_to_wrap.gamelogic.setWord\[17\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3650_ net254 vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
X_3581_ net276 vssd1 vssd1 vccd1 vccd1 _0113_ sky130_fd_sc_hd__inv_2
X_2601_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[5\] _1275_ _1285_ team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2532_ net472 team_10_WB.instance_to_wrap.buffer.temp_guess\[4\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4202_ clknet_leaf_12_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[64\]
+ _0191_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[64\] sky130_fd_sc_hd__dfrtp_1
X_2463_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] net197 team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\]
+ _1191_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2394_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _1089_ _1158_ net575 vssd1
+ vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4133_ clknet_leaf_9_wb_clk_i _0604_ _0132_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ clknet_leaf_21_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[1\]
+ _0084_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3015_ team_10_WB.instance_to_wrap.gamelogic.setWord\[4\] net190 vssd1 vssd1 vccd1
+ vccd1 _1502_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2491__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout246_A net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3917_ net247 vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__inv_2
X_3848_ net241 vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3779_ net271 vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout201_X net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout121 net124 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
Xfanout110 net115 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__buf_2
XFILLER_0_11_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout132 _1183_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_2
Xfanout165 net166 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input6_X net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 net145 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
X_4532__344 vssd1 vssd1 vccd1 vccd1 _4532__344/HI net344 sky130_fd_sc_hd__conb_1
Xfanout187 _0994_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
Xfanout176 _1440_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
Xfanout198 _0826_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4041__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4191__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2473__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1963_ team_10_WB.instance_to_wrap.gamelogic.setWord\[31\] _0874_ _0877_ net157 vssd1
+ vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4682_ net182 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1894_ team_10_WB.instance_to_wrap.host_col\[3\] vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__inv_2
X_3702_ net235 vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3633_ net252 vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3564_ net290 vssd1 vssd1 vccd1 vccd1 _0096_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1953__B net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3495_ net250 vssd1 vssd1 vccd1 vccd1 _0027_ sky130_fd_sc_hd__inv_2
X_2515_ net224 _1225_ net193 vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o21ai_1
X_4516__328 vssd1 vssd1 vccd1 vccd1 _4516__328/HI net328 sky130_fd_sc_hd__conb_1
X_2446_ _1187_ _1196_ net584 net129 vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__o2bb2a_1
X_4116_ clknet_leaf_9_wb_clk_i _0587_ _0115_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[51\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2377_ _1126_ _1129_ _1128_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__a21oi_1
X_4047_ clknet_leaf_14_wb_clk_i _0532_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4207__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3008__A2 net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4603__378 vssd1 vssd1 vccd1 vccd1 _4603__378/HI net378 sky130_fd_sc_hd__conb_1
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1990__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4064__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2455__B1 _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4407__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1966__C1 net157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1981__A2 net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _1666_ _1667_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__nor2_1
X_2300_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[7\] _1076_ _1077_
+ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__and3_1
X_2231_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] _0803_ vssd1 vssd1 vccd1
+ vccd1 _1013_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3333__X _1713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2162_ _0942_ _0944_ _0956_ net642 vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a22o_1
X_2093_ team_10_WB.instance_to_wrap.dispFSM.guesses\[19\] net113 net140 net641 vssd1
+ vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_42 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_642 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2995_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[33\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[34\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[35\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[36\]
+ net161 vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__a41o_1
XFILLER_0_12_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4087__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3410__A2 _1703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1946_ _0845_ _0855_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__nand2_1
X_4665_ net431 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[4] sky130_fd_sc_hd__buf_2
X_1877_ net215 vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
X_4596_ net200 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3616_ net251 vssd1 vssd1 vccd1 vccd1 _0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3547_ net290 vssd1 vssd1 vccd1 vccd1 _0079_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3478_ team_10_WB.instance_to_wrap.host_row2\[47\] net174 _1708_ team_10_WB.instance_to_wrap.host_row1\[79\]
+ _1850_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__a221o_1
XANTENNA__2795__A net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2429_ net511 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[39\]
+ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__a22o_1
XANTENNA__3477__A2 net173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3403__B _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2437__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2988__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1874__A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1963__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4538__350 vssd1 vssd1 vccd1 vccd1 _4538__350/HI net350 sky130_fd_sc_hd__conb_1
XFILLER_0_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input41_A wbs_dat_i[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3468__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2780_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _1390_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold207 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[43\] vssd1 vssd1 vccd1
+ vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
X_4450_ clknet_leaf_27_wb_clk_i net502 _0433_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold229 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[38\] vssd1 vssd1 vccd1
+ vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ net174 net171 net181 vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__or3_1
Xhold218 team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\] vssd1 vssd1 vccd1 vccd1
+ net675 sky130_fd_sc_hd__dlygate4sd3_1
X_4381_ clknet_leaf_2_wb_clk_i _0766_ _0364_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[18\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__3947__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3332_ team_10_WB.instance_to_wrap.host_row1\[72\] _1708_ _1711_ net304 _1706_ vssd1
+ vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3263_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] _1653_ net514 vssd1 vssd1
+ vccd1 vccd1 _1656_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3459__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3194_ _1390_ _1611_ _1614_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and3b_1
X_2214_ net12 net11 net14 net13 vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__or4_2
XFILLER_0_56_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2145_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\] team_10_WB.instance_to_wrap.gamelogic.rights\[0\]
+ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__or2_1
X_2076_ team_10_WB.instance_to_wrap.dispFSM.guesses\[36\] net109 net135 net698 vssd1
+ vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__o22a_1
XANTENNA__3947__Q team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_A _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_344 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2978_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[20\] net160 _1488_ net214
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[20\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3395__B2 team_10_WB.instance_to_wrap.host_row2\[67\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1929_ net226 _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__nor2_1
X_4648_ net417 vssd1 vssd1 vccd1 vccd1 la_data_out[18] sky130_fd_sc_hd__buf_2
XFILLER_0_60_946 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_136 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4579_ net199 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4102__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3083__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4609__384 vssd1 vssd1 vccd1 vccd1 _4609__384/HI net384 sky130_fd_sc_hd__conb_1
XFILLER_0_35_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1875__Y _0800_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3138__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2212__B net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2897__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4616__388 vssd1 vssd1 vccd1 vccd1 _4616__388/HI net388 sky130_fd_sc_hd__conb_1
Xhold90 team_10_WB.instance_to_wrap.keypadFSMPlayer.prev_key\[5\] vssd1 vssd1 vccd1
+ vccd1 net547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3074__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3950_ clknet_leaf_22_wb_clk_i _0013_ net284 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.keypadFSMPlayer.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2901_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[14\] net155 net122 net608
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[6\]
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_34_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3881_ net276 vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__inv_2
X_2832_ _1405_ _1433_ _1434_ _1432_ vssd1 vssd1 vccd1 vccd1 _0001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2763_ _1379_ _1380_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[22\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4502_ net314 vssd1 vssd1 vccd1 vccd1 ADR_O[9] sky130_fd_sc_hd__buf_2
XFILLER_0_53_261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_935 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2694_ net600 _1009_ _1339_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[1\]
+ sky130_fd_sc_hd__o21bai_1
X_4433_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[30\]
+ _0416_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4125__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4364_ clknet_leaf_2_wb_clk_i _0749_ _0347_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_3315_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[1\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\]
+ _1682_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__and3_1
X_4295_ clknet_leaf_15_wb_clk_i _0685_ _0284_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2018__C_N net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3246_ _1608_ _1645_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__or2_1
XANTENNA__4275__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3177_ _1283_ _1599_ _1601_ net195 vssd1 vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2128_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] team_10_WB.instance_to_wrap.buffer.temp_guess\[5\]
+ _0926_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3065__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2059_ net569 net143 net107 net594 vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1056 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_932 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2040__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2207__B _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4148__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2223__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4298__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[19] sky130_fd_sc_hd__clkbuf_4
X_3100_ net207 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\] net191 _1544_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[86\] sky130_fd_sc_hd__a31o_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 gpio_out[35] sky130_fd_sc_hd__buf_2
X_4080_ clknet_leaf_13_wb_clk_i _0551_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3031_ team_10_WB.instance_to_wrap.gamelogic.setWord\[12\] team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[12\]
+ net188 vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__mux2_1
XANTENNA__2893__A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3933_ net237 vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__inv_2
X_3864_ net261 vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__inv_2
X_2815_ _0514_ _0515_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3795_ net272 vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2746_ team_10_WB.instance_to_wrap.clock_div.count\[17\] _1367_ vssd1 vssd1 vccd1
+ vccd1 _1369_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2133__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2677_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] _1327_ _1318_ vssd1
+ vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4416_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[13\]
+ _0399_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4347_ clknet_leaf_19_wb_clk_i _0737_ _0336_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[70\]
+ sky130_fd_sc_hd__dfstp_1
X_4278_ clknet_leaf_17_wb_clk_i _0668_ _0267_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[1\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_fanout181_X net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3229_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\]
+ _1632_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[16\] vssd1 vssd1 vccd1 vccd1
+ _1636_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_38_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2261__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[38\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4440__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3580_ net263 vssd1 vssd1 vccd1 vccd1 _0112_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2600_ _1270_ _1284_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2531_ net467 team_10_WB.instance_to_wrap.buffer.temp_guess\[5\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_286 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4201_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[63\]
+ _0190_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[63\] sky130_fd_sc_hd__dfrtp_1
X_2462_ net474 net131 _1204_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2393_ team_10_WB.instance_to_wrap.keypadFSMHost.unlocked _1093_ _1158_ net550 vssd1
+ vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__a22o_1
X_4132_ clknet_leaf_9_wb_clk_i _0603_ _0131_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[67\]
+ sky130_fd_sc_hd__dfrtp_1
X_4063_ clknet_leaf_21_wb_clk_i team_10_WB.instance_to_wrap.uart_transmitter.next_state\[0\]
+ _0083_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3014_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[3\] net185 _1501_ net206
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[43\] sky130_fd_sc_hd__o211a_1
XFILLER_0_64_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4313__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4629__398 vssd1 vssd1 vccd1 vccd1 _4629__398/HI net398 sky130_fd_sc_hd__conb_1
XFILLER_0_59_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3916_ net264 vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout239_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3847_ net259 vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__inv_2
XANTENNA__4463__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ net283 vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__inv_2
X_2729_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ _1358_ _1177_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_14_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout122 net124 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout133 _1183_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_2
Xfanout155 _1182_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_2
Xfanout188 net189 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__clkbuf_2
Xfanout177 net178 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout199 net201 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_2
Xfanout166 _0872_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1877__A net215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_26_wb_clk_i_X clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__2473__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1962_ team_10_WB.instance_to_wrap.gamelogic.setWord\[23\] net147 vssd1 vssd1 vccd1
+ vccd1 _0877_ sky130_fd_sc_hd__or2_1
X_4681_ net435 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[20] sky130_fd_sc_hd__buf_2
X_1893_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[0\] vssd1 vssd1 vccd1 vccd1
+ _0817_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3701_ net235 vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__inv_2
XANTENNA__1984__B1 net119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3632_ net252 vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3563_ net289 vssd1 vssd1 vccd1 vccd1 _0095_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3066__X team_10_WB.instance_to_wrap.hostdisp.nextBottom\[69\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2514_ _1226_ _1229_ net193 vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__and3b_1
X_3494_ net254 vssd1 vssd1 vccd1 vccd1 _0026_ sky130_fd_sc_hd__inv_2
X_4555__367 vssd1 vssd1 vccd1 vccd1 _4555__367/HI net367 sky130_fd_sc_hd__conb_1
X_2445_ _0836_ net194 vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4115_ clknet_leaf_9_wb_clk_i _0586_ _0114_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[50\]
+ sky130_fd_sc_hd__dfrtp_1
X_2376_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] _1084_ _1148_
+ _1149_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout189_A _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4046_ clknet_leaf_14_wb_clk_i _0531_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3413__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4223__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[85\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4209__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_58_Left_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4359__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3404__B1 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _0822_ team_10_WB.instance_to_wrap.gamelogic.state\[1\] team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ _0988_ team_10_WB.instance_to_wrap.gamelogic.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _1012_ sky130_fd_sc_hd__a311o_1
X_2161_ _0942_ _0943_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__a21o_1
X_2092_ team_10_WB.instance_to_wrap.dispFSM.guesses\[20\] net109 net136 net701 vssd1
+ vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2446__B2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2994_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[37\] net158 vssd1 vssd1 vccd1
+ vccd1 _1493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _0845_ _0855_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4664_ net184 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1876_ net214 vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ net199 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_1
X_3615_ net252 vssd1 vssd1 vccd1 vccd1 _0147_ sky130_fd_sc_hd__inv_2
X_3546_ net286 vssd1 vssd1 vccd1 vccd1 _0078_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3477_ team_10_WB.instance_to_wrap.host_row2\[87\] net173 net180 team_10_WB.instance_to_wrap.host_row2\[63\]
+ net304 vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__a221o_1
XANTENNA__2134__A0 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2428_ net192 _1185_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2_1
X_2359_ _1124_ _1134_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__xnor2_1
X_4029_ clknet_leaf_11_wb_clk_i _0514_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_4644__413 vssd1 vssd1 vccd1 vccd1 _4644__413/HI net413 sky130_fd_sc_hd__conb_1
XFILLER_0_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4031__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_657 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_156 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4181__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input34_A wbs_adr_i[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[25\] vssd1 vssd1 vccd1
+ vccd1 net665 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3328__Y _1708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold219 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[17\] vssd1 vssd1 vccd1
+ vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
X_4380_ clknet_leaf_7_wb_clk_i _0765_ _0363_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[17\]
+ sky130_fd_sc_hd__dfstp_2
X_3400_ _1686_ _1698_ _1776_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__or3_1
XANTENNA__2903__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3331_ team_10_WB.instance_to_wrap.host_row2\[56\] net180 net167 team_10_WB.instance_to_wrap.host_row2\[72\]
+ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3262_ net629 _1653_ _1655_ vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__o21a_1
X_2213_ net39 net38 net10 net9 vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3193_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\] vssd1 vssd1 vccd1 vccd1 _1614_
+ sky130_fd_sc_hd__a21o_1
X_2144_ team_10_WB.instance_to_wrap.gamelogic.incorrect\[2\] team_10_WB.instance_to_wrap.gamelogic.incorrect\[1\]
+ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__a21o_1
X_2075_ net565 net143 net107 net576 vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__a22o_1
XANTENNA__4054__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3092__A1 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2977_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[19\] net164 _1488_ team_10_WB.instance_to_wrap.gamelogic.letter\[3\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[19\]
+ sky130_fd_sc_hd__o22a_1
XANTENNA__3395__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ team_10_WB.instance_to_wrap.host_col\[3\] net225 vssd1 vssd1 vccd1 vccd1 _0851_
+ sky130_fd_sc_hd__or2_2
X_4647_ net416 vssd1 vssd1 vccd1 vccd1 la_data_out[17] sky130_fd_sc_hd__buf_2
XFILLER_0_60_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4578_ net199 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_1
X_3529_ net271 vssd1 vssd1 vccd1 vccd1 _0061_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_wb_clk_i clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3386__A2 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_52_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold91 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[13\] vssd1 vssd1 vccd1 vccd1
+ net548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[17\] vssd1 vssd1 vccd1 vccd1
+ net537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4077__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2900_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[13\] net156 net125 net494
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[5\]
+ sky130_fd_sc_hd__a22o_1
X_3880_ net261 vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
X_2831_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3377__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2762_ team_10_WB.instance_to_wrap.clock_div.count\[21\] team_10_WB.instance_to_wrap.clock_div.count\[20\]
+ team_10_WB.instance_to_wrap.clock_div.count\[22\] _1374_ vssd1 vssd1 vccd1 vccd1
+ _1380_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4501_ net313 vssd1 vssd1 vccd1 vccd1 ADR_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2693_ _1009_ _1238_ _1339_ _1340_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_transmitter.next_state\[0\]
+ sky130_fd_sc_hd__a22o_1
X_4432_ clknet_leaf_26_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[29\]
+ _0415_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4363_ clknet_leaf_2_wb_clk_i _0748_ _0346_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_3314_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\] team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__nand2_2
X_4294_ clknet_leaf_17_wb_clk_i _0684_ _0283_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[17\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3245_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[2\] vssd1 vssd1 vccd1 vccd1 _1645_
+ sky130_fd_sc_hd__a21oi_1
X_3176_ _1582_ _1600_ _0906_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2127_ _0919_ _0928_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout269_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2058_ team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] net111 net139 net639 vssd1
+ vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_538 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_944 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3368__A2 net177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3359__A2 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2567__B1 team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[1] sky130_fd_sc_hd__clkbuf_4
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 gpio_out[36] sky130_fd_sc_hd__buf_2
X_3030_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] _1509_ net206 vssd1 vssd1
+ vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[51\] sky130_fd_sc_hd__mux2_1
XANTENNA__2893__B net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_321 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3932_ net265 vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3863_ net275 vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__inv_2
X_2814_ _1413_ _1418_ _1416_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__a21o_1
X_3794_ net281 vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2745_ _1367_ _1368_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[16\]
+ sky130_fd_sc_hd__nor2_1
X_2676_ _1318_ _1328_ _1329_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[5\]
+ sky130_fd_sc_hd__and3_1
X_4415_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[12\]
+ _0398_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2420__Y _1182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1972__B net147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout304 net6 vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__buf_4
X_4346_ clknet_leaf_18_wb_clk_i net583 _0335_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[69\]
+ sky130_fd_sc_hd__dfrtp_1
X_4277_ clknet_leaf_14_wb_clk_i _0667_ _0266_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4392__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3228_ net644 _1633_ _1635_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__o21a_1
XANTENNA__2089__A2 net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_X net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _1586_ _1587_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_473 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4115__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2234__A team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4222__Q team_10_WB.instance_to_wrap.host_row2\[84\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2530_ net462 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\] _1233_ vssd1 vssd1
+ vccd1 vccd1 _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2461_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[5\] net208 team_10_WB.instance_to_wrap.hostdisp.curr_word\[21\]
+ _1189_ net129 vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__o221a_1
X_4200_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[62\]
+ _0189_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[62\] sky130_fd_sc_hd__dfrtp_1
X_2392_ net2 net596 _1158_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4131_ clknet_leaf_2_wb_clk_i _0602_ _0130_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[66\]
+ sky130_fd_sc_hd__dfrtp_1
X_4062_ clknet_leaf_14_wb_clk_i net513 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_3013_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] net190 vssd1 vssd1 vccd1
+ vccd1 _1501_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3915_ net247 vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3440__B2 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3846_ net242 vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_390 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3777_ net292 vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout301_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2728_ team_10_WB.instance_to_wrap.clock_div.count\[10\] _1356_ vssd1 vssd1 vccd1
+ vccd1 _1358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2951__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2659_ _1310_ _1317_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout112 net115 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_2
X_4329_ clknet_leaf_17_wb_clk_i _0719_ _0318_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[52\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout134 _0919_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_2
Xfanout145 _0912_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
Xfanout156 _1181_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_4
Xfanout178 _1399_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
Xfanout167 _1710_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_4
Xfanout189 _0994_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_4
XANTENNA__4138__CLK clknet_leaf_10_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4288__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2942__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2473__A2 net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1961_ team_10_WB.instance_to_wrap.gamelogic.setWord\[24\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[32\]
+ vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__o22a_1
XANTENNA__3422__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ net236 vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ net182 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_1
X_1892_ team_10_WB.instance_to_wrap.lcdPlayer.currentState\[0\] vssd1 vssd1 vccd1
+ vccd1 _0816_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1984__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[14\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1984__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3631_ net253 vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3562_ net289 vssd1 vssd1 vccd1 vccd1 _0094_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2933__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2513_ net224 _1225_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] vssd1
+ vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3493_ net251 vssd1 vssd1 vccd1 vccd1 _0025_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2444_ net581 net133 _1185_ _1195_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2375_ team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] _1075_ _1141_
+ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__a21o_1
X_4114_ clknet_leaf_9_wb_clk_i _0585_ _0113_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__2161__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4045_ clknet_leaf_14_wb_clk_i _0530_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2449__C1 _1190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2139__A net134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2464__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4566__442 vssd1 vssd1 vccd1 vccd1 net442 _4566__442/LO sky130_fd_sc_hd__conb_1
XANTENNA__4430__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout137_X net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3829_ net249 vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2924__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_555 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2455__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1966__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[29\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3608__A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2915__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4303__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4453__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2160_ _0936_ _0941_ _0954_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__a21o_1
X_4589__453 vssd1 vssd1 vccd1 vccd1 net453 _4589__453/LO sky130_fd_sc_hd__conb_1
X_2091_ team_10_WB.instance_to_wrap.dispFSM.guesses\[29\] net143 net108 net597 vssd1
+ vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2993_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\] net158 _1492_ net212
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[31\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_452 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1944_ _0858_ _0866_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4522__334 vssd1 vssd1 vccd1 vccd1 _4522__334/HI net334 sky130_fd_sc_hd__conb_1
X_4663_ net184 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3614_ net251 vssd1 vssd1 vccd1 vccd1 _0146_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1875_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1 vccd1
+ _0800_ sky130_fd_sc_hd__inv_2
XANTENNA__2906__B1 net121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4594_ net199 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3545_ net286 vssd1 vssd1 vccd1 vccd1 _0077_ sky130_fd_sc_hd__inv_2
X_3476_ team_10_WB.instance_to_wrap.host_row1\[55\] _1699_ net169 team_10_WB.instance_to_wrap.host_row1\[63\]
+ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__a22o_1
X_2427_ net185 _1186_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nor2_1
XANTENNA__3331__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2358_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1133_ _1132_ _1117_
+ _1100_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__o2111a_1
X_2289_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__inv_2
X_4028_ clknet_leaf_11_wb_clk_i _0513_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.currentState\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2437__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3970__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4326__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4476__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input27_A wbs_adr_i[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4506__318 vssd1 vssd1 vccd1 vccd1 _4506__318/HI net318 sky130_fd_sc_hd__conb_1
XFILLER_0_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3389__B1 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold209 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\] vssd1 vssd1 vccd1 vccd1
+ net666 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3330_ _1683_ _1687_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3261_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[8\] _1653_ net296 vssd1 vssd1
+ vccd1 vccd1 _1655_ sky130_fd_sc_hd__a21oi_1
X_2212_ net19 net8 net33 net30 vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__or4_1
X_3192_ _1389_ _1611_ _1613_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2143_ team_10_WB.instance_to_wrap.correct\[1\] team_10_WB.instance_to_wrap.correct\[0\]
+ team_10_WB.instance_to_wrap.correct\[2\] vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__o21a_1
XANTENNA__3993__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2074_ team_10_WB.instance_to_wrap.dispFSM.guesses\[38\] net111 net138 net692 vssd1
+ vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2976_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[18\] net160 _1488_ net216
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[18\]
+ sky130_fd_sc_hd__o22a_1
X_1927_ net229 _0848_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4646_ net415 vssd1 vssd1 vccd1 vccd1 la_data_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_fanout214_A team_10_WB.instance_to_wrap.gamelogic.letter\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4577_ net199 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3528_ net246 vssd1 vssd1 vccd1 vccd1 _0060_ sky130_fd_sc_hd__inv_2
X_3459_ team_10_WB.instance_to_wrap.dispFSM.guesses\[62\] _1701_ _1717_ team_10_WB.instance_to_wrap.dispFSM.guesses\[6\]
+ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_680 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2997__A team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[4\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2897__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold81 team_10_WB.instance_to_wrap.host_row1\[43\] vssd1 vssd1 vccd1 vccd1 net538
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 team_10_WB.instance_to_wrap.keypadFSMPlayer.unlocked vssd1 vssd1 vccd1 vccd1
+ net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 team_10_WB.instance_to_wrap.uart_transmitter.clk_count\[7\] vssd1 vssd1 vccd1
+ vccd1 net527 sky130_fd_sc_hd__dlygate4sd3_1
X_2830_ _1430_ _1431_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3339__Y _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2761_ team_10_WB.instance_to_wrap.clock_div.count\[22\] _1378_ vssd1 vssd1 vccd1
+ vccd1 _1379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4500_ net312 vssd1 vssd1 vccd1 vccd1 ADR_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_5_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2692_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] _1241_ vssd1 vssd1
+ vccd1 vccd1 _1340_ sky130_fd_sc_hd__or2_1
XANTENNA_1 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4431_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[28\]
+ _0414_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_13_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4362_ clknet_leaf_12_wb_clk_i _0747_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_4293_ clknet_leaf_14_wb_clk_i _0683_ _0282_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[16\]
+ sky130_fd_sc_hd__dfstp_1
X_3313_ net210 _1686_ _1688_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\]
+ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__and4b_4
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3244_ _1610_ _1644_ net298 vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__a21oi_1
X_3175_ _0887_ _0894_ _0891_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3531__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2126_ net213 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0928_ sky130_fd_sc_hd__mux2_1
XANTENNA__4171__CLK clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout164_A net166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2057_ team_10_WB.instance_to_wrap.dispFSM.guesses\[63\] net144 net108 net627 vssd1
+ vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__a22o_1
X_4528__340 vssd1 vssd1 vccd1 vccd1 _4528__340/HI net340 sky130_fd_sc_hd__conb_1
XFILLER_0_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_422 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2959_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[1\] _1480_ _1481_ vssd1
+ vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_X net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4629_ net398 vssd1 vssd1 vccd1 vccd1 irq[2] sky130_fd_sc_hd__buf_2
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3706__A net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_809 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2223__C net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4044__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[21] sky130_fd_sc_hd__clkbuf_4
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4194__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4018__RESET_B net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3931_ net248 vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__inv_2
X_3862_ net261 vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
X_2813_ _1415_ _1417_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__or2_1
X_3793_ net292 vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2744_ team_10_WB.instance_to_wrap.clock_div.count\[16\] _1365_ _1177_ vssd1 vssd1
+ vccd1 vccd1 _1368_ sky130_fd_sc_hd__o21ai_1
X_2675_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[3\]
+ _1321_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\] vssd1 vssd1 vccd1
+ vccd1 _1329_ sky130_fd_sc_hd__a31o_1
X_4414_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[11\]
+ _0397_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2430__A _0993_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4345_ clknet_leaf_16_wb_clk_i _0735_ _0334_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[68\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4276_ clknet_leaf_1_wb_clk_i _0666_ _0265_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3227_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[15\] _1633_ _1612_ vssd1
+ vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__a21oi_1
XANTENNA__2494__B1 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ _1560_ _1585_ _1584_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ team_10_WB.instance_to_wrap.dispFSM.guesses\[3\] net115 net136 team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] net197 vssd1 vssd1 vccd1
+ vccd1 _1539_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_X net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2485__B1 _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1897__Y _0821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_wb_clk_i clknet_2_3__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_X clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2460_ net486 _1184_ _1203_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4130_ clknet_leaf_10_wb_clk_i _0601_ _0129_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[65\]
+ sky130_fd_sc_hd__dfrtp_1
X_2391_ net526 _1158_ _1159_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4061_ clknet_leaf_15_wb_clk_i _0546_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3012_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[2\] net185 _1500_ net203
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[42\] sky130_fd_sc_hd__o211a_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3914_ net243 vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2425__A net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3845_ net248 vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3776_ net293 vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout127_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2431__Y _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2727_ _1180_ _1355_ _1357_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[9\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_15_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2951__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[3\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2658_ _1222_ _1234_ _1225_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o21bai_2
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_2
XFILLER_0_1_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2589_ _1272_ _1273_ _0902_ _0908_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__o2bb2a_1
Xfanout146 net147 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_4
Xfanout124 _1473_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
Xfanout135 net137 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
X_4328_ clknet_leaf_16_wb_clk_i _0718_ _0317_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[51\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout179 _1727_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_4
Xfanout168 _1710_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_2
X_4259_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[2\]
+ _0248_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_input1_A gpio_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _0873_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_42_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1993__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2942__A1 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3407__C1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ team_10_WB.instance_to_wrap.gamelogic.setWord\[25\] net146 net116 team_10_WB.instance_to_wrap.gamelogic.setWord\[33\]
+ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_16_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1891_ team_10_WB.instance_to_wrap.lcdPlayer.nextState\[3\] vssd1 vssd1 vccd1 vccd1
+ _0815_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1984__A2 net149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4382__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ net267 vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3561_ net289 vssd1 vssd1 vccd1 vccd1 _0093_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2512_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] _1226_ _1228_ vssd1
+ vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3492_ net250 vssd1 vssd1 vccd1 vccd1 _0024_ sky130_fd_sc_hd__inv_2
X_2443_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net185 vssd1 vssd1 vccd1
+ vccd1 _1195_ sky130_fd_sc_hd__or2_1
X_2374_ _0871_ _1147_ _1087_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__a21oi_1
X_4113_ clknet_leaf_10_wb_clk_i _0584_ _0112_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_4044_ clknet_leaf_14_wb_clk_i _0529_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2449__B1 _1191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4408__Q team_10_WB.instance_to_wrap.hostdisp.curr_word\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2426__Y _1187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3413__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout244_A net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3828_ net264 vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3759_ net280 vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__inv_2
XANTENNA__4105__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_567 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input4_X net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4255__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2215__D _1000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1966__A2 _0874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2090_ team_10_WB.instance_to_wrap.dispFSM.guesses\[22\] net111 net139 net690 vssd1
+ vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2527__X _1233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[30\] net161 _1491_ team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[30\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1943_ _0844_ net196 vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__and2_1
X_4662_ net182 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_1
X_4561__373 vssd1 vssd1 vccd1 vccd1 _4561__373/HI net373 sky130_fd_sc_hd__conb_1
XFILLER_0_43_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1874_ net213 vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3613_ net251 vssd1 vssd1 vccd1 vccd1 _0145_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4593_ net200 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2422__B _1181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4128__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3544_ net284 vssd1 vssd1 vccd1 vccd1 _0076_ sky130_fd_sc_hd__inv_2
X_3475_ team_10_WB.instance_to_wrap.host_row1\[47\] _1693_ _1703_ team_10_WB.instance_to_wrap.host_row1\[71\]
+ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2426_ _0993_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__nor2_2
XANTENNA__4278__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout194_A _0991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2357_ _0823_ _0828_ _1859_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__and3_1
X_2288_ team_10_WB.instance_to_wrap.host_col\[3\] net226 team_10_WB.instance_to_wrap.host_col\[0\]
+ net225 vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__or4b_2
X_4027_ clknet_leaf_1_wb_clk_i net466 _0074_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_895 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4545__357 vssd1 vssd1 vccd1 vccd1 _4545__357/HI net357 sky130_fd_sc_hd__conb_1
XFILLER_0_38_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3619__A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4420__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3260_ net475 _1651_ _1654_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o21a_1
X_2211_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__or4_1
X_3191_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__or2_1
X_2142_ _0916_ _0935_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__or2_1
X_2073_ net558 net144 net108 net589 vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__a22o_1
XANTENNA__3092__A3 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[17\] net164 _1488_ net217
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[17\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1926_ net229 _0848_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nor2_1
X_4645_ net414 vssd1 vssd1 vccd1 vccd1 la_data_out[15] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Left_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout207_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4576_ net199 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3527_ net246 vssd1 vssd1 vccd1 vccd1 _0059_ sky130_fd_sc_hd__inv_2
X_3458_ team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] net168 _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[14\]
+ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3389_ team_10_WB.instance_to_wrap.dispFSM.guesses\[59\] _1701_ net181 team_10_WB.instance_to_wrap.dispFSM.guesses\[35\]
+ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__a22o_1
X_2409_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[3\] team_10_WB.instance_to_wrap.clock_div.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout197_X net197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3068__A0 team_10_WB.instance_to_wrap.gamelogic.setWord\[22\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_228 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4443__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3174__A team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[15\] vssd1 vssd1 vccd1 vccd1
+ net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 team_10_WB.instance_to_wrap.host_row1\[76\] vssd1 vssd1 vccd1 vccd1 net539
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 team_10_WB.instance_to_wrap.host_row1\[53\] vssd1 vssd1 vccd1 vccd1 net528
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 team_10_WB.instance_to_wrap.keypadFSMHost.prev_key\[3\] vssd1 vssd1 vccd1
+ vccd1 net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2760_ _1377_ _1378_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[21\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2034__B2 team_10_WB.instance_to_wrap.dispFSM.msg\[6\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2691_ team_10_WB.instance_to_wrap.uart_transmitter.state\[0\] _1246_ _1238_ vssd1
+ vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__a21oi_1
XANTENNA_2 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[27\]
+ _0413_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_35_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4634__403 vssd1 vssd1 vccd1 vccd1 _4634__403/HI net403 sky130_fd_sc_hd__conb_1
X_4361_ clknet_leaf_12_wb_clk_i _0004_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2742__C1 _1177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3312_ _1691_ _1692_ net282 vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a21oi_1
X_4292_ clknet_leaf_19_wb_clk_i net578 _0281_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_3243_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[1\] team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[0\]
+ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3960__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3174_ team_10_WB.instance_to_wrap.dispFSM.msg\[6\] _1550_ vssd1 vssd1 vccd1 vccd1
+ _1599_ sky130_fd_sc_hd__or2_1
XANTENNA__3023__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4316__CLK clknet_leaf_18_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2125_ _0919_ _0927_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__and2_1
XANTENNA__2428__A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2056_ team_10_WB.instance_to_wrap.dispFSM.guesses\[56\] net113 net140 net638 vssd1
+ vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout157_A _0873_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__B1 _1717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4466__CLK clknet_leaf_1_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2958_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\] _0832_ net163 vssd1 vssd1 vccd1
+ vccd1 _1481_ sky130_fd_sc_hd__a41o_1
XFILLER_0_8_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_434 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1909_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\] vssd1 vssd1 vccd1 vccd1
+ _0832_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4628_ net397 vssd1 vssd1 vccd1 vccd1 irq[1] sky130_fd_sc_hd__buf_2
XANTENNA__4151__Q net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2889_ team_10_WB.instance_to_wrap.buffer.Rx_byte\[6\] net1 _1469_ vssd1 vssd1 vccd1
+ vccd1 _1470_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4559_ net371 vssd1 vssd1 vccd1 vccd1 SEL_O[1] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_9_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3722__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3461__B1 _1719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2801__A net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput50 net50 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[23] sky130_fd_sc_hd__clkbuf_4
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA_input42_X net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4489__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3930_ net242 vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3452__B1 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3861_ net262 vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__inv_2
X_2812_ _0816_ _0817_ net177 vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__mux2_1
X_3792_ net293 vssd1 vssd1 vccd1 vccd1 _0324_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2743_ team_10_WB.instance_to_wrap.clock_div.count\[15\] team_10_WB.instance_to_wrap.clock_div.count\[16\]
+ _1364_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2674_ _1327_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__inv_2
X_4413_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[10\]
+ _0396_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__2430__B _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4344_ clknet_leaf_18_wb_clk_i _0734_ _0333_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[67\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_1_375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload11_A clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4275_ clknet_leaf_1_wb_clk_i _0665_ _0264_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_3226_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1632_ _1634_ vssd1
+ vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout274_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3157_ _1560_ _1584_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2108_ team_10_WB.instance_to_wrap.dispFSM.guesses\[4\] net114 net141 team_10_WB.instance_to_wrap.dispFSM.guesses\[12\]
+ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ net204 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[40\] net187 _1538_
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[80\] sky130_fd_sc_hd__a31o_1
X_2039_ team_10_WB.instance_to_wrap.dispFSM.guesses\[73\] net110 net137 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__o22a_1
XANTENNA__3443__B1 net167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Left_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2237__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[6\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2237__B2 team_10_WB.instance_to_wrap.gamelogic.setWord\[0\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4011__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4161__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_952 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2390_ _0858_ _1158_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__nor2_1
X_4060_ clknet_leaf_15_wb_clk_i _0545_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3011_ team_10_WB.instance_to_wrap.gamelogic.setWord\[2\] net192 vssd1 vssd1 vccd1
+ vccd1 _1500_ sky130_fd_sc_hd__or2_1
XANTENNA__3425__B1 _1693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3913_ net257 vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__inv_2
XANTENNA__2425__B _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3844_ net260 vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3775_ net280 vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3537__A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2726_ _1356_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2657_ _1222_ _1225_ _1227_ _1234_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[2\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2588_ _0898_ _0901_ _0907_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__and3_1
Xfanout114 net115 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_2
Xfanout136 net137 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_2
X_4327_ clknet_leaf_16_wb_clk_i _0717_ _0316_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[50\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout147 net150 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
Xfanout125 _1472_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout169 _1704_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_4
X_4258_ clknet_leaf_3_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[1\]
+ _0247_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout158 net159 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
X_3209_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[8\] _1621_ _1623_ vssd1 vssd1
+ vccd1 vccd1 _0535_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4189_ clknet_leaf_8_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[51\]
+ _0178_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[51\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__3416__B1 _1720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4034__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4184__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2942__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_0_Left_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold190 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[34\] vssd1 vssd1 vccd1
+ vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1969__B1 net117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1890_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_20ms\[5\] vssd1 vssd1 vccd1 vccd1
+ _0814_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3560_ net289 vssd1 vssd1 vccd1 vccd1 _0092_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2511_ _1225_ _1227_ _1222_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3491_ net253 vssd1 vssd1 vccd1 vccd1 _0023_ sky130_fd_sc_hd__inv_2
X_2442_ net505 net131 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[31\]
+ vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__a22o_1
XANTENNA__3343__C1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2373_ _1137_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__or2_1
X_4112_ clknet_leaf_2_wb_clk_i _0583_ _0111_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_4043_ clknet_leaf_13_wb_clk_i _0528_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4057__CLK clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3827_ net254 vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3758_ net296 vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2709_ _1345_ _1346_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2924__A2 net156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3689_ net236 vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2128__A0 team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_45_Left_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2256__A team_10_WB.instance_to_wrap.gamelogic.setWord\[33\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2991_ net631 net158 _1492_ team_10_WB.instance_to_wrap.gamelogic.letter\[5\] vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[29\] sky130_fd_sc_hd__a22o_1
XFILLER_0_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1942_ _0819_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__nand2_1
X_4661_ net430 vssd1 vssd1 vccd1 vccd1 la_data_out[31] sky130_fd_sc_hd__buf_2
X_1873_ team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1 vccd1 vccd1
+ _0798_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3612_ net280 vssd1 vssd1 vccd1 vccd1 _0144_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4592_ net456 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XANTENNA__2906__A2 net153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3374__X _1752_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clknet_2_0__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3543_ net290 vssd1 vssd1 vccd1 vccd1 _0075_ sky130_fd_sc_hd__inv_2
XANTENNA__3815__A net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3474_ team_10_WB.instance_to_wrap.dispFSM.guesses\[31\] net171 net168 team_10_WB.instance_to_wrap.dispFSM.guesses\[55\]
+ _1846_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__a221o_1
X_2425_ net197 _0942_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clknet_0_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3331__A2 net180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2356_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] _1119_ vssd1 vssd1 vccd1
+ vccd1 _1132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout187_A _0994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2287_ _1064_ _1063_ team_10_WB.instance_to_wrap.gamelogic.rights\[0\] vssd1 vssd1
+ vccd1 vccd1 _0644_ sky130_fd_sc_hd__mux2_1
X_4026_ clknet_leaf_1_wb_clk_i net463 _0073_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4154__Q net71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3725__A net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_25_wb_clk_i_X clknet_leaf_25_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4372__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3389__A2 _1701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2210_ _0806_ _0996_ net194 _0945_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__a2bb2o_1
X_3190_ net478 net172 vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__nor2_1
X_2141_ _0916_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__nor2_1
X_2072_ team_10_WB.instance_to_wrap.dispFSM.guesses\[40\] net113 net140 net658 vssd1
+ vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2974_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[16\] net160 _1488_ team_10_WB.instance_to_wrap.gamelogic.letter\[0\]
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[16\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_wb_clk_i clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1925_ net2 net3 net300 vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2052__A2 net115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4644_ net413 vssd1 vssd1 vccd1 vccd1 la_data_out[14] sky130_fd_sc_hd__buf_2
XANTENNA__3001__B2 team_10_WB.instance_to_wrap.gamelogic.letter\[2\] vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
X_4575_ net199 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3526_ net246 vssd1 vssd1 vccd1 vccd1 _0058_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4395__CLK clknet_leaf_6_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3457_ team_10_WB.instance_to_wrap.host_row1\[78\] _1708_ _1829_ _1830_ vssd1 vssd1
+ vccd1 vccd1 _1831_ sky130_fd_sc_hd__a211o_1
XANTENNA__4149__Q net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3388_ team_10_WB.instance_to_wrap.dispFSM.guesses\[75\] _1715_ _1720_ team_10_WB.instance_to_wrap.dispFSM.guesses\[11\]
+ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__a221o_1
X_2408_ _1164_ _1167_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_4_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2339_ _1110_ _1111_ _1113_ _1114_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4009_ clknet_leaf_21_wb_clk_i _0497_ net285 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4512__324 vssd1 vssd1 vccd1 vccd1 _4512__324/HI net324 sky130_fd_sc_hd__conb_1
Xhold50 team_10_WB.instance_to_wrap.host_row1\[55\] vssd1 vssd1 vccd1 vccd1 net507
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input32_A wbs_adr_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 team_10_WB.instance_to_wrap.host_row1\[46\] vssd1 vssd1 vccd1 vccd1 net518
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 team_10_WB.instance_to_wrap.host_row1\[44\] vssd1 vssd1 vccd1 vccd1 net529
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 team_10_WB.instance_to_wrap.host_row1\[49\] vssd1 vssd1 vccd1 vccd1 net540
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_2_1__f_wb_clk_i_X clknet_2_1__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 team_10_WB.instance_to_wrap.host_row1\[51\] vssd1 vssd1 vccd1 vccd1 net551
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4118__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4268__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2253__B net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2690_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[10\] _1336_ _1338_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_3 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ clknet_leaf_12_wb_clk_i _0003_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.nextState\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3311_ net178 net489 vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4291_ clknet_leaf_19_wb_clk_i _0681_ _0280_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[14\]
+ sky130_fd_sc_hd__dfstp_1
X_3242_ net503 _1610_ net298 vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__a21oi_1
X_3173_ _0903_ _1298_ _1598_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__a21o_1
X_2124_ net212 team_10_WB.instance_to_wrap.buffer.temp_guess\[7\] _0926_ vssd1 vssd1
+ vccd1 vccd1 _0927_ sky130_fd_sc_hd__mux2_1
XANTENNA__2428__B _1185_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2055_ team_10_WB.instance_to_wrap.dispFSM.guesses\[57\] net110 net135 net710 vssd1
+ vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2957_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[11\] team_10_WB.instance_to_wrap.hostdisp.curr_word\[12\]
+ team_10_WB.instance_to_wrap.hostdisp.curr_word\[14\] _0833_ net163 vssd1 vssd1 vccd1
+ vccd1 _1480_ sky130_fd_sc_hd__a41o_1
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1908_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[7\] vssd1 vssd1 vccd1 vccd1
+ _0831_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2888_ net224 team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\]
+ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__and3b_1
X_4627_ net396 vssd1 vssd1 vccd1 vccd1 irq[0] sky130_fd_sc_hd__buf_2
XFILLER_0_60_725 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2981__A0 net212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4558_ net370 vssd1 vssd1 vccd1 vccd1 SEL_O[0] sky130_fd_sc_hd__buf_2
XFILLER_0_60_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4489_ clknet_leaf_7_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[46\]
+ _0472_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[46\]
+ sky130_fd_sc_hd__dfstp_1
X_3509_ net250 vssd1 vssd1 vccd1 vccd1 _0041_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4410__CLK clknet_leaf_2_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_777 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4657__426 vssd1 vssd1 vccd1 vccd1 _4657__426/HI net426 sky130_fd_sc_hd__conb_1
Xoutput51 net51 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 gpio_oeb[35] sky130_fd_sc_hd__buf_2
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3860_ net263 vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2811_ _1413_ _1415_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3791_ net281 vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2742_ team_10_WB.instance_to_wrap.clock_div.count\[15\] _1364_ _1366_ _1177_ vssd1
+ vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.next_count\[15\] sky130_fd_sc_hd__o211a_1
XFILLER_0_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4412_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[9\]
+ _0395_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[9\]
+ sky130_fd_sc_hd__dfstp_1
X_2673_ team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] team_10_WB.instance_to_wrap.uart_receiver.clk_count\[5\]
+ _1324_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__and3_1
X_4343_ clknet_leaf_16_wb_clk_i _0733_ _0332_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[66\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_10_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4274_ clknet_leaf_1_wb_clk_i _0664_ _0263_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3225_ _1612_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__nor2_1
XANTENNA__3034__S net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2494__A2 net130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4433__CLK clknet_leaf_9_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3156_ _1569_ _1574_ _1573_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3087_ _0790_ net204 vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2107_ team_10_WB.instance_to_wrap.dispFSM.guesses\[13\] net143 net107 net484 vssd1
+ vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__a22o_1
X_2038_ team_10_WB.instance_to_wrap.dispFSM.guesses\[74\] net112 net139 team_10_WB.instance_to_wrap.dispFSM.msg\[2\]
+ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3989_ clknet_leaf_29_wb_clk_i team_10_WB.instance_to_wrap.clock_div.next_count\[26\]
+ _0057_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.clock_div.count\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2954__B1 _1478_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_316 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3950__CLK clknet_leaf_22_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1996__A1 team_10_WB.instance_to_wrap.gamelogic.setWord\[5\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4306__CLK clknet_leaf_19_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4518__330 vssd1 vssd1 vccd1 vccd1 _4518__330/HI net330 sky130_fd_sc_hd__conb_1
XANTENNA__3370__B1 net174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output63_A net201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4456__CLK clknet_leaf_27_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3010_ team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[1\] net186 _1499_ net207
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.nextBottom\[41\] sky130_fd_sc_hd__o211a_1
XFILLER_0_64_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3912_ net240 vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__inv_2
X_3843_ net247 vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4605__380 vssd1 vssd1 vccd1 vccd1 _4605__380/HI net380 sky130_fd_sc_hd__conb_1
X_3774_ net295 vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3029__S net190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2725_ team_10_WB.instance_to_wrap.clock_div.count\[7\] team_10_WB.instance_to_wrap.clock_div.count\[8\]
+ team_10_WB.instance_to_wrap.clock_div.count\[9\] _1351_ vssd1 vssd1 vccd1 vccd1
+ _1356_ sky130_fd_sc_hd__and4_2
X_2656_ _1307_ _1316_ _1314_ _1228_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_state\[1\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3361__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2164__A1 _0942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2587_ net5 _0902_ _0904_ _1271_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2217__D_N net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4326_ clknet_leaf_17_wb_clk_i _0716_ _0315_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[49\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout126 _1191_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_4
Xfanout115 _0913_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout137 _0914_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_2
Xfanout148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
Xfanout159 _0873_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__buf_2
X_4257_ clknet_leaf_0_wb_clk_i team_10_WB.instance_to_wrap.gamelogic.nextState\[0\]
+ _0246_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3208_ net172 _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__nor2_1
X_4188_ clknet_leaf_2_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.nextBottom\[50\]
+ _0177_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row2\[50\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__2467__A2 net129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3139_ _1286_ _1554_ _1565_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_59_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3973__CLK clknet_leaf_28_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4582__450 vssd1 vssd1 vccd1 vccd1 net450 _4582__450/LO sky130_fd_sc_hd__conb_1
XFILLER_0_64_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4329__CLK clknet_leaf_17_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2927__B1 net120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_566 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3352__B1 _1715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 team_10_WB.instance_to_wrap.dispFSM.guesses\[54\] vssd1 vssd1 vccd1 vccd1
+ net637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[30\] vssd1 vssd1 vccd1
+ vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3407__A1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output101_A net184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2918__B1 net125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2510_ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[2\] team_10_WB.instance_to_wrap.uart_receiver.bit_index\[1\]
+ team_10_WB.instance_to_wrap.uart_receiver.bit_index\[0\] vssd1 vssd1 vccd1 vccd1
+ _1227_ sky130_fd_sc_hd__and3_1
X_3490_ net267 vssd1 vssd1 vccd1 vccd1 _0022_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clknet_2_2__leaf_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2441_ net531 net130 net127 team_10_WB.instance_to_wrap.hostdisp.curr_word\[32\]
+ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__a22o_1
XANTENNA__3343__B1 _1704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2372_ _1131_ _1135_ _1096_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__a21oi_1
X_4111_ clknet_leaf_7_wb_clk_i _0582_ _0110_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.host_row1\[46\]
+ sky130_fd_sc_hd__dfrtp_1
X_4042_ clknet_leaf_13_wb_clk_i _0527_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__2449__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3996__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_305 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3826_ net258 vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2909__B1 net122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_15_wb_clk_i_X clknet_leaf_15_wb_clk_i vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3757_ net285 vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2708_ team_10_WB.instance_to_wrap.clock_div.count\[1\] team_10_WB.instance_to_wrap.clock_div.count\[0\]
+ team_10_WB.instance_to_wrap.clock_div.count\[2\] vssd1 vssd1 vccd1 vccd1 _1346_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__2385__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[0\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3688_ net237 vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__inv_2
X_4573__449 vssd1 vssd1 vccd1 vccd1 net449 _4573__449/LO sky130_fd_sc_hd__conb_1
X_2639_ _0946_ _1304_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.nextState\[0\]
+ sky130_fd_sc_hd__nand2_1
X_4309_ clknet_leaf_12_wb_clk_i _0699_ _0298_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[32\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4001__CLK clknet_leaf_24_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4151__CLK clknet_leaf_11_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3022__C1 net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2376__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[2\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3325__B1 net169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3480__X _1853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__2256__B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2990_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[28\] net161 _1491_ net214
+ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[28\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1941_ net229 _0848_ _0851_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4660_ net429 vssd1 vssd1 vccd1 vccd1 la_data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1872_ team_10_WB.instance_to_wrap.gamelogic.setWord\[3\] vssd1 vssd1 vccd1 vccd1
+ _0797_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3087__B net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3611_ net254 vssd1 vssd1 vccd1 vccd1 _0143_ sky130_fd_sc_hd__inv_2
X_4591_ net455 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XANTENNA__2367__A1 team_10_WB.instance_to_wrap.host_message_reg.setLetter\[4\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3542_ net237 vssd1 vssd1 vccd1 vccd1 _0074_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3473_ team_10_WB.instance_to_wrap.dispFSM.msg\[7\] net169 _1844_ _1845_ vssd1 vssd1
+ vccd1 vccd1 _1846_ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_7 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2424_ net197 _0942_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__nor2_4
X_2355_ _1128_ _1129_ _1126_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__a21bo_1
X_2286_ _0940_ _1064_ _1065_ _1063_ team_10_WB.instance_to_wrap.gamelogic.rights\[1\]
+ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4174__CLK clknet_leaf_26_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4025_ clknet_leaf_1_wb_clk_i net468 _0072_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.buffer.temp_guess\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4662__A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3809_ net292 vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_812 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4170__Q team_10_WB.instance_to_wrap.host_message_reg.setLetter\[3\] vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_X net302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4618__390 vssd1 vssd1 vccd1 vccd1 _4618__390/HI net390 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_54_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3188__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3010__A2 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4047__CLK clknet_leaf_14_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4197__CLK clknet_leaf_8_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2140_ _0822_ net218 vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand2_1
X_2071_ team_10_WB.instance_to_wrap.dispFSM.guesses\[41\] net109 net135 net715 vssd1
+ vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2037__B1 net137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1045 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_2973_ team_10_WB.instance_to_wrap.gamelogic.indexCorrect\[2\] net126 _1486_ _1487_
+ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__nand4_4
XFILLER_0_57_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1924_ net300 net3 vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ net412 vssd1 vssd1 vccd1 vccd1 la_data_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_60_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4574_ net201 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_1
X_3525_ net245 vssd1 vssd1 vccd1 vccd1 _0057_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3037__S net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3456_ team_10_WB.instance_to_wrap.host_row1\[46\] _1693_ net174 team_10_WB.instance_to_wrap.host_row2\[46\]
+ _1826_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout297_A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_3387_ team_10_WB.instance_to_wrap.dispFSM.guesses\[51\] net168 _1719_ team_10_WB.instance_to_wrap.dispFSM.guesses\[67\]
+ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__a22o_1
X_2407_ _1168_ _1169_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2338_ _0811_ _1093_ _1107_ _1108_ _1109_ vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2269_ team_10_WB.instance_to_wrap.gamelogic.setWord\[30\] net213 vssd1 vssd1 vccd1
+ vccd1 _1051_ sky130_fd_sc_hd__nand2_1
X_4008_ clknet_leaf_19_wb_clk_i _0496_ net285 vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.msg\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_19_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Left_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4551__363 vssd1 vssd1 vccd1 vccd1 _4551__363/HI net363 sky130_fd_sc_hd__conb_1
Xhold40 team_10_WB.instance_to_wrap.message_reg.msg\[2\] vssd1 vssd1 vccd1 vccd1 net497
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[6\] vssd1 vssd1 vccd1
+ vccd1 net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 team_10_WB.instance_to_wrap.message_reg.msg\[3\] vssd1 vssd1 vccd1 vccd1 net530
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input25_A wbs_adr_i[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold51 team_10_WB.instance_to_wrap.dispFSM.guesses\[7\] vssd1 vssd1 vccd1 vccd1 net508
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 team_10_WB.instance_to_wrap.host_row1\[54\] vssd1 vssd1 vccd1 vccd1 net552
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 team_10_WB.instance_to_wrap.uart_receiver.clk_count\[4\] vssd1 vssd1 vccd1
+ vccd1 net541 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2518__C net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2990__B2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3310_ _1684_ _1689_ _1690_ net177 vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__or4b_1
XFILLER_0_46_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4290_ clknet_leaf_18_wb_clk_i net563 _0279_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3241_ net512 _1642_ _1643_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__o21a_1
X_3172_ _1290_ _1597_ team_10_WB.instance_to_wrap.dispFSM.msg\[5\] vssd1 vssd1 vccd1
+ vccd1 _1598_ sky130_fd_sc_hd__o21a_1
X_2123_ _0918_ _0925_ _0922_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__a21oi_4
X_2054_ team_10_WB.instance_to_wrap.dispFSM.guesses\[58\] net111 net138 net657 vssd1
+ vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4212__CLK clknet_leaf_3_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3470__A2 net175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2956_ team_10_WB.instance_to_wrap.hostdisp.curr_word\[13\] net158 vssd1 vssd1 vccd1
+ vccd1 _1479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1907_ team_10_WB.instance_to_wrap.keypadFSMHost.state\[5\] vssd1 vssd1 vccd1 vccd1
+ _0830_ sky130_fd_sc_hd__inv_2
X_2887_ net193 _1468_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.temp_byte\[5\]
+ sky130_fd_sc_hd__and2_1
X_4626_ net395 vssd1 vssd1 vccd1 vccd1 gpio_out[37] sky130_fd_sc_hd__buf_2
XFILLER_0_60_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4362__CLK clknet_leaf_12_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout212_A team_10_WB.instance_to_wrap.gamelogic.letter\[7\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4494__306 vssd1 vssd1 vccd1 vccd1 _4494__306/HI net306 sky130_fd_sc_hd__conb_1
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4557_ net369 vssd1 vssd1 vccd1 vccd1 DAT_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_12_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3508_ net246 vssd1 vssd1 vccd1 vccd1 _0040_ sky130_fd_sc_hd__inv_2
X_4488_ clknet_leaf_1_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_guesses\[45\]
+ _0471_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_guesses\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4535__347 vssd1 vssd1 vccd1 vccd1 _4535__347/HI net347 sky130_fd_sc_hd__conb_1
XANTENNA__3291__A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3439_ team_10_WB.instance_to_wrap.host_row2\[101\] team_10_WB.instance_to_wrap.dispFSM.guesses\[5\]
+ net303 vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__mux2_1
XANTENNA__2249__B1 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3461__A2 net181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput52 net52 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
Xoutput63 net201 vssd1 vssd1 vccd1 vccd1 gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 wbs_dat_o[26] sky130_fd_sc_hd__clkbuf_4
XANTENNA__2488__B1 net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input28_X net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_804 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__4235__CLK clknet_leaf_21_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3452__A2 _1699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4182__D team_10_WB.instance_to_wrap.hostdisp.nextBottom\[44\] vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4385__CLK clknet_leaf_7_wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2810_ _1415_ vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ net296 vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_222 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2741_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__inv_2
XANTENNA__2963__B2 net216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__3095__B net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4411_ clknet_leaf_9_wb_clk_i team_10_WB.instance_to_wrap.hostdisp.next_curr_word\[8\]
+ _0394_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.hostdisp.curr_word\[8\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2672_ net541 _1324_ _1326_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.uart_receiver.next_clk_count\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4342_ clknet_leaf_17_wb_clk_i _0732_ _0331_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.dispFSM.guesses\[65\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_2_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_4273_ clknet_leaf_0_wb_clk_i _0663_ _0262_ vssd1 vssd1 vccd1 vccd1 team_10_WB.instance_to_wrap.gamelogic.letter\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_3224_ team_10_WB.instance_to_wrap.lcdPlayer.cnt_500hz\[14\] _1632_ vssd1 vssd1 vccd1
+ vccd1 _1633_ sky130_fd_sc_hd__and2_1
.ends

